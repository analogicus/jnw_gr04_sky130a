magic
tech sky130A
magscale 1 2
timestamp 1744580037
<< locali >>
rect -3056 22216 -2744 22328
rect -1600 22280 -1360 22720
rect -1026 21404 -834 22396
rect 9922 20906 10002 21080
rect 2244 19985 3868 20177
rect 2244 18475 2436 19985
rect 8770 19230 8830 19458
rect 7370 19170 8830 19230
rect 2244 18469 2558 18475
rect 2244 18421 2504 18469
rect 2552 18421 2558 18469
rect 2244 18415 2558 18421
rect -2949 14305 -841 15625
rect 2244 15164 2436 18415
rect 4920 18224 5348 18416
rect 5156 18026 5348 18224
rect 7370 18230 7430 19170
rect 7370 18229 8830 18230
rect 7370 18223 8944 18229
rect 7370 18221 8890 18223
rect 7363 18175 8890 18221
rect 8938 18175 8944 18223
rect 7363 18170 8944 18175
rect 7363 18154 7427 18170
rect 8766 18169 8944 18170
rect 7363 18102 7369 18154
rect 7421 18102 7427 18154
rect 7363 18096 7427 18102
rect 5156 17870 5174 18026
rect 5330 17870 5348 18026
rect 5156 17392 5348 17870
rect 8884 17481 8944 17625
rect 4645 17195 4821 17356
rect 5011 17200 5348 17392
rect 4645 17031 4651 17195
rect 4815 17031 4821 17195
rect 4645 17025 4821 17031
rect 5165 17064 5664 17124
rect 5165 16276 5225 17064
rect 5852 16786 5984 16846
rect 8084 16055 8144 16181
rect 5471 16007 8144 16055
rect 5411 15995 8144 16007
rect 2244 14972 9032 15164
rect 2244 12667 2436 14972
rect 8840 12667 9032 14972
rect 126 12475 9032 12667
<< viali >>
rect 4898 22772 5062 22936
rect -5278 22522 -5122 22678
rect -3596 22480 -3368 22720
rect -2514 22486 -2286 22714
rect 9922 21080 10002 21148
rect 7990 20918 8070 20986
rect 2504 18421 2552 18469
rect 1967 16599 2147 16779
rect 8890 18175 8938 18223
rect 7369 18102 7421 18154
rect 5174 17870 5330 18026
rect 8884 17625 8944 17673
rect 4651 17031 4815 17195
rect 5804 16786 5852 16846
rect 5411 16007 5471 16055
<< metal1 >>
rect 5290 22942 5466 22948
rect 4886 22936 5290 22942
rect -2754 22877 -2514 22883
rect -2754 22813 4400 22877
rect -3602 22720 -3362 22732
rect -2754 22720 -2514 22813
rect -5284 22678 -5116 22690
rect -5284 22522 -5278 22678
rect -5122 22522 -5116 22678
rect -5284 22084 -5116 22522
rect -3602 22480 -3596 22720
rect -3368 22714 -2274 22720
rect -3368 22486 -2514 22714
rect -2286 22486 -2274 22714
rect 4336 22640 4400 22813
rect 4886 22772 4898 22936
rect 5062 22772 5290 22936
rect 4886 22766 5290 22772
rect 5290 22760 5466 22766
rect 4330 22576 4336 22640
rect 4400 22576 4406 22640
rect -3368 22480 -2274 22486
rect -3602 22468 -3362 22480
rect -5284 21916 -4716 22084
rect -4884 20271 -4716 21916
rect -1518 21919 972 22111
rect 2028 21919 2808 22111
rect -1518 21335 -1326 21919
rect 4440 21883 4446 21947
rect 4510 21883 4516 21947
rect 1268 21461 1332 21467
rect 4468 21461 4532 21467
rect 1184 21257 1190 21449
rect 1268 21391 1332 21397
rect 1382 21257 1388 21449
rect 2362 21397 2368 21461
rect 2432 21397 2438 21461
rect -1621 20561 -450 20753
rect 2368 20432 2432 21397
rect 4468 21391 4532 21397
rect 8138 21302 8314 21308
rect 7272 21126 8138 21302
rect 7990 20992 8070 21126
rect 8138 21120 8314 21126
rect 9722 21074 9728 21154
rect 9808 21148 10014 21154
rect 9808 21080 9922 21148
rect 10002 21080 10014 21148
rect 9808 21074 10014 21080
rect 7978 20986 8082 20992
rect 7978 20918 7990 20986
rect 8070 20918 8082 20986
rect 7978 20912 8082 20918
rect 2368 20368 2632 20432
rect 2568 19832 2632 20368
rect 2568 19768 3032 19832
rect 2968 18896 3032 19768
rect 2968 18832 3482 18896
rect 2968 18762 3032 18768
rect 2660 18475 2720 18481
rect 2492 18469 2660 18475
rect 2492 18421 2504 18469
rect 2552 18421 2660 18469
rect 2492 18415 2660 18421
rect 2660 18409 2720 18415
rect 2967 18267 3027 18273
rect 2967 18176 3027 18207
rect 3418 18117 3482 18832
rect 8884 18223 8944 18235
rect 8884 18175 8890 18223
rect 8938 18175 8944 18223
rect 7363 18160 7427 18166
rect 4968 18154 7427 18160
rect 3418 18053 3858 18117
rect 4968 18102 7369 18154
rect 7421 18102 7427 18154
rect 4968 18096 7427 18102
rect 7363 18090 7427 18096
rect 3788 17776 3852 18053
rect 4864 18026 5342 18032
rect 4864 17870 5174 18026
rect 5330 17870 5342 18026
rect 4864 17864 5342 17870
rect 3775 17584 4504 17776
rect 5470 17621 6384 17681
rect 8884 17679 8944 18175
rect 8872 17673 8956 17679
rect 8872 17625 8884 17673
rect 8944 17625 8956 17673
rect 4925 17201 5101 17207
rect 4639 17195 4925 17201
rect 4639 17031 4651 17195
rect 4815 17031 4925 17195
rect 4639 17025 4925 17031
rect 4925 17019 5101 17025
rect 5470 17022 5530 17621
rect 8872 17619 8956 17625
rect 5470 16956 5530 16962
rect 5798 16846 5858 16858
rect 5418 16786 5804 16846
rect 5852 16786 5858 16846
rect 1955 16779 3913 16785
rect 1955 16599 1967 16779
rect 2147 16661 3913 16779
rect 4167 16661 4343 16667
rect 2147 16599 4167 16661
rect 1955 16593 4167 16599
rect 3747 16485 4167 16593
rect 4167 16479 4343 16485
rect 5418 16127 5478 16786
rect 5798 16774 5858 16786
rect 5411 16061 5478 16127
rect 5399 16055 5483 16061
rect 5399 16007 5411 16055
rect 5471 16007 5483 16055
rect 5399 16001 5483 16007
<< via1 >>
rect 5290 22766 5466 22942
rect 4336 22576 4400 22640
rect 4446 21883 4510 21947
rect 1268 21397 1332 21461
rect 2368 21397 2432 21461
rect 4468 21397 4532 21461
rect 8138 21126 8314 21302
rect 9728 21074 9808 21154
rect 2968 18768 3032 18832
rect 2660 18415 2720 18475
rect 2967 18207 3027 18267
rect 4925 17025 5101 17201
rect 5470 16962 5530 17022
rect 4167 16485 4343 16661
<< metal2 >>
rect 5284 22766 5290 22942
rect 5466 22937 9346 22942
rect 5466 22771 9175 22937
rect 9341 22771 9350 22937
rect 5466 22766 9346 22771
rect 4336 22640 4400 22646
rect 4336 21947 4400 22576
rect 4446 21947 4510 21953
rect 4336 21883 4446 21947
rect 4446 21877 4510 21883
rect 2368 21461 2432 21467
rect 1262 21397 1268 21461
rect 1332 21397 2368 21461
rect 2432 21397 4468 21461
rect 4532 21397 4538 21461
rect 2368 21391 2432 21397
rect 8635 21302 8801 21306
rect 8132 21126 8138 21302
rect 8314 21297 8806 21302
rect 8314 21131 8635 21297
rect 8801 21131 8806 21297
rect 9728 21154 9808 21160
rect 8314 21126 8806 21131
rect 8635 21122 8801 21126
rect 9573 21074 9582 21154
rect 9652 21074 9728 21154
rect 9728 21068 9808 21074
rect 2962 18768 2968 18832
rect 3032 18768 3038 18832
rect 2968 18579 3032 18768
rect 2968 18514 3032 18523
rect 2654 18415 2660 18475
rect 2720 18415 2726 18475
rect 2660 18362 2720 18415
rect 2653 18306 2662 18362
rect 2718 18306 2727 18362
rect 2967 18354 3027 18363
rect 2660 18304 2720 18306
rect 2967 18267 3027 18298
rect 2961 18207 2967 18267
rect 3027 18207 3033 18267
rect 5240 17201 5406 17205
rect 4919 17025 4925 17201
rect 5101 17196 5411 17201
rect 5101 17030 5240 17196
rect 5406 17030 5411 17196
rect 5101 17025 5411 17030
rect 5240 17021 5406 17025
rect 5464 16962 5470 17022
rect 5530 16962 5536 17022
rect 5470 16818 5530 16962
rect 5470 16753 5530 16762
rect 4463 16661 4629 16665
rect 4161 16485 4167 16661
rect 4343 16656 4634 16661
rect 4343 16490 4463 16656
rect 4629 16490 4634 16656
rect 4343 16485 4634 16490
rect 4463 16481 4629 16485
<< via2 >>
rect 9175 22771 9341 22937
rect 8635 21131 8801 21297
rect 9582 21074 9652 21154
rect 2968 18523 3032 18579
rect 2662 18306 2718 18362
rect 2967 18298 3027 18354
rect 5240 17030 5406 17196
rect 5470 16762 5530 16818
rect 4463 16490 4629 16656
<< metal3 >>
rect 9170 22937 9346 22942
rect 9170 22771 9175 22937
rect 9341 22771 9346 22937
rect 8630 21297 8806 21302
rect 8630 21131 8635 21297
rect 8801 21131 8806 21297
rect 8630 20772 8806 21131
rect 9170 21154 9346 22771
rect 9577 21154 9657 21159
rect 9170 21074 9582 21154
rect 9652 21074 9657 21154
rect 9170 20772 9346 21074
rect 9577 21069 9657 21074
rect 2963 18579 3037 18584
rect 2963 18523 2968 18579
rect 3032 18523 3037 18579
rect 2963 18518 3037 18523
rect 2657 18362 2723 18367
rect 2657 18306 2662 18362
rect 2718 18306 2723 18362
rect 2968 18359 3032 18518
rect 2657 18301 2723 18306
rect 2962 18354 3032 18359
rect 2660 18162 2720 18301
rect 2962 18298 2967 18354
rect 3027 18298 3032 18354
rect 2962 18293 3032 18298
rect 2652 18098 2658 18162
rect 2722 18098 2728 18162
rect 2968 17925 3032 18293
rect 5235 17196 5730 17201
rect 5235 17030 5240 17196
rect 5406 17030 5730 17196
rect 9342 17034 9992 17201
rect 5235 17025 5730 17030
rect 9218 17025 9992 17034
rect 5465 16818 5535 16823
rect 5465 16762 5470 16818
rect 5530 16762 5535 16818
rect 5465 16757 5535 16762
rect 5470 16661 5530 16757
rect 4458 16656 5730 16661
rect 4458 16490 4463 16656
rect 4629 16490 5730 16656
rect 4458 16485 5730 16490
rect 9218 16485 10118 16661
<< via3 >>
rect 2658 18098 2722 18162
<< metal4 >>
rect 2657 18162 2723 18163
rect 2657 18098 2658 18162
rect 2722 18098 2723 18162
rect 2657 18097 2723 18098
rect 2660 17919 2720 18097
use JNWTR_RPPO8  x3 ../JNW_TR_SKY130A
timestamp 1744566163
transform -1 0 -2956 0 -1 25640
box 0 0 2744 3440
use JNWTR_RPPO4  x4 ../JNW_TR_SKY130A
timestamp 1744227008
transform -1 0 -996 0 -1 25638
box 0 0 1880 3440
use JNWTR_DFRNQNX1_CV  x6 ../JNW_TR_SKY130A
timestamp 1744566163
transform 0 -1 9390 -1 0 17831
box -150 -120 2130 3960
use JNWTR_SCX1_CV  x9 ../JNW_TR_SKY130A
timestamp 1744580037
transform 1 0 8005 0 -1 20946
box -150 -120 2130 1720
use JNWTR_CAPX1  xc1 ../JNW_TR_SKY130A
timestamp 1737500400
transform -1 0 3614 0 -1 17955
box 0 0 1080 1080
use PTAT  xp1 ../JNW_GR04_SKY130A
timestamp 1744566163
transform -1 0 -6307 0 1 14265
box -5108 -265 5202 7780
use Current_mirror  xp2 ../JNW_GR04_SKY130A
timestamp 1744566163
transform -1 0 2054 0 1 12793
box -204 -524 3168 9318
use Opamp_test  xp3 ../JNW_GR04_SKY130A
timestamp 1744566163
transform 0 -1 9056 1 0 16153
box 2222 1594 6906 6420
use JNWATR_NCH_2C1F2  xr1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 -1 5072 -1 0 18320
box -184 -128 1208 928
<< labels >>
flabel locali 5165 16276 5225 16336 0 FreeSans 1600 0 0 0 OUT
port 2 nsew
flabel metal3 9809 16485 9985 16661 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel metal3 9816 17025 9992 17201 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 14697 25807
<< end >>
