*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR04_lpe.spi
#else
.include ../../../work/xsch/JNW_GR04.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.save i(Vbias)
.save i(R1)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control

set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 1u 0



foreach vtemp -40 -20 0 20 40 80 125

  option temp=$vtemp
  tran 1n 100n

  set fend = .raw
  write {cicname}_$vtemp$fend
end

quit

.endc

.end
