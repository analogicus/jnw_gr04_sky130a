magic
tech sky130A
magscale 1 2
timestamp 1744495200
<< checkpaint >>
rect -368934881474191040 -368934881474191040 -184467440737095520 4826
use pnp_05v5 xb1 ../sky130_fd_pr
transform 1 0 0 0 1 0
box 0 0 -368934881474191040 -368934881474191040
use pnp_05v5 xb2 ../sky130_fd_pr
transform 1 0 0 0 1 -368934881474191040
box 0 -368934881474191040 -368934881474191040 -737869762948382080
use JNWTR_CAPX1 xc1 ../JNW_TR_SKY130A
transform 1 0 -368934881474191040 0 1 0
box -368934881474191040 0 -368934881474189975 1080
use JNWATR_PCH_4C5F0 xm1 ../JNW_ATR_SKY130A
transform 1 0 -368934881474189952 0 1 0
box -368934881474189952 0 -368934881474188805 800
use JNWATR_PCH_4C5F0 xm2 ../JNW_ATR_SKY130A
transform 1 0 -368934881474189952 0 1 800
box -368934881474189952 800 -368934881474188805 1600
use JNWATR_PCH_4C5F0 xm3 ../JNW_ATR_SKY130A
transform 1 0 -368934881474189952 0 1 1600
box -368934881474189952 1600 -368934881474188805 2400
use Opamp_test xo1 ../JNW_GR04_SKY130A
transform 1 0 -368934881474188800 0 1 0
box -368934881474188800 0 -368934881474184622 4826
use JNWTR_RPPO16 xr1 ../JNW_TR_SKY130A
transform 1 0 -368934881474184640 0 1 0
box -368934881474184640 0 -368934881474180175 3440
<< labels >>
<< properties >>
string FIXED_BBOX -368934881474191040 -368934881474191040 -184467440737095520 4826
<< end >>
