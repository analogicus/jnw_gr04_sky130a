magic
tech sky130A
timestamp 1744367994
<< locali >>
rect 2110 2904 2206 3235
rect 2686 3123 2833 3133
rect 2686 3045 2716 3123
rect 2794 3045 2833 3123
rect 2686 2880 2833 3045
rect 2110 2612 2206 2661
rect 1317 2364 1437 2609
rect 1987 2556 2206 2612
rect 2110 2251 2206 2556
rect 2686 2649 2806 2680
rect 2686 2237 2833 2649
rect 3313 2264 3409 2656
rect 2713 2225 2833 2237
rect 2110 1744 2206 2001
rect 3313 1697 3409 1976
rect 2110 896 2206 1074
rect 2686 896 2833 1098
rect 3313 896 3409 1074
rect 2110 893 3409 896
rect 2110 803 2497 893
rect 2587 803 2932 893
rect 3022 803 3409 893
rect 2110 800 3409 803
<< viali >>
rect 2716 3045 2794 3123
rect 1759 2382 1849 2472
rect 2497 803 2587 893
rect 2932 803 3022 893
<< metal1 >>
rect 2496 3126 2580 3243
rect 2941 3126 3025 3131
rect 2496 3123 3025 3126
rect 2496 3045 2716 3123
rect 2794 3045 3025 3123
rect 2496 3042 3025 3045
rect 2496 2876 2580 3042
rect 2941 2876 3025 3042
rect 2302 2532 2398 2727
rect 2622 2532 2654 2648
rect 2865 2532 2897 2632
rect 2301 2500 2897 2532
rect 2302 2475 2398 2500
rect 1753 2472 2398 2475
rect 1753 2382 1759 2472
rect 1849 2382 2398 2472
rect 3121 2467 3217 2696
rect 2504 2466 3217 2467
rect 1753 2379 2398 2382
rect 2500 2383 3217 2466
rect 2500 2221 2584 2383
rect 2931 2315 3025 2383
rect 2929 2221 3025 2315
rect 2302 1857 2398 2029
rect 2622 1895 2654 1977
rect 2865 1893 2897 1977
rect 2302 1825 2897 1857
rect 2302 1667 2398 1825
rect 2622 1743 2654 1825
rect 2865 1745 2897 1825
rect 3121 1629 3217 2068
rect 2302 1282 2398 1544
rect 2494 1180 2590 1592
rect 2622 1343 2654 1447
rect 2865 1369 2897 1489
rect 2865 1321 2897 1366
rect 2929 1183 3025 1562
rect 3121 1242 3217 1513
rect 2494 893 2590 1150
rect 2494 803 2497 893
rect 2587 803 2590 893
rect 2494 797 2590 803
rect 2929 893 3025 1150
rect 2929 803 2932 893
rect 3022 803 3025 893
rect 2929 797 3025 803
use JNWTR_RPPO4  x2 ../JNW_TR_SKY130A
timestamp 1744227008
transform -1 0 2051 0 1 904
box 0 0 940 1720
use JNWATR_PCH_4C1F2  xb1 ../JNW_ATR_SKY130A
timestamp 1744227008
transform -1 0 2734 0 1 2580
box -92 -64 668 464
use JNWATR_PCH_4C1F2  xb2
timestamp 1744227008
transform 1 0 2785 0 1 2580
box -92 -64 668 464
use JNWATR_PCH_4C1F2  xi1
timestamp 1744227008
transform -1 0 2734 0 1 1925
box -92 -64 668 464
use JNWATR_PCH_4C1F2  xi2
timestamp 1744227008
transform 1 0 2785 0 1 1925
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xm1_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform -1 0 2734 0 1 998
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xm1_1
timestamp 1734044400
transform -1 0 2734 0 1 1397
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xm2_0
timestamp 1734044400
transform 1 0 2785 0 1 998
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xm2_1
timestamp 1734044400
transform 1 0 2785 0 1 1397
box -92 -64 668 464
<< labels >>
flabel metal1 2865 1893 2897 1977 0 FreeSans 800 0 0 0 VIN
port 2 nsew
flabel metal1 2622 1895 2654 1977 0 FreeSans 800 0 0 0 VIP
port 4 nsew
flabel locali 2110 2904 2206 3235 0 FreeSans 800 0 0 0 VSS
port 6 nsew
flabel metal1 2496 2876 2580 3238 0 FreeSans 800 0 0 0 VDD
port 8 nsew
flabel metal1 3121 1629 3217 2068 0 FreeSans 800 0 0 0 Vo
port 10 nsew
<< end >>
