magic
tech sky130A
timestamp 1744566163
<< locali >>
rect -48 4441 149 4537
rect 239 4441 621 4537
rect -48 4309 48 4441
rect 525 4357 621 4441
rect 868 -51 964 82
rect 868 -139 1063 -51
rect 1441 -51 1537 38
rect 1153 -139 1537 -51
rect 868 -147 1537 -139
<< viali >>
rect 149 4441 239 4537
rect 1063 -139 1153 -49
<< metal1 >>
rect -102 4563 637 4659
rect 144 4543 240 4563
rect 144 4537 242 4543
rect 144 4441 149 4537
rect 239 4441 242 4537
rect 144 4435 242 4441
rect 706 4436 1347 4532
rect 80 4084 112 4087
rect 80 3941 112 4067
rect 80 3680 112 3683
rect 80 3645 112 3648
rect 77 3520 80 3552
rect 112 3520 115 3552
rect 80 3274 112 3277
rect 80 3239 112 3242
rect 77 3123 80 3155
rect 112 3123 115 3155
rect 80 2873 112 2876
rect 80 2838 112 2841
rect 77 2731 80 2763
rect 112 2731 115 2763
rect 80 2471 112 2474
rect 80 2436 112 2439
rect 77 2307 80 2339
rect 112 2307 115 2339
rect 80 2070 112 2073
rect 80 2035 112 2038
rect 77 1927 80 1959
rect 112 1927 115 1959
rect 80 1677 112 1680
rect 80 1642 112 1645
rect 77 1515 80 1547
rect 112 1515 115 1547
rect 80 1277 112 1280
rect 80 1242 112 1245
rect 77 1097 80 1129
rect 112 1097 115 1129
rect 80 876 112 879
rect 80 841 112 844
rect 77 717 80 749
rect 112 717 115 749
rect 80 476 112 479
rect 80 441 112 444
rect 77 322 80 354
rect 112 322 115 354
rect 77 78 80 110
rect 112 78 115 110
rect 144 12 240 4435
rect 336 4219 488 4315
rect 706 3917 802 4436
rect 996 4062 1028 4065
rect 996 4027 1028 4030
rect 336 3821 819 3917
rect 993 3905 996 3937
rect 1028 3905 1031 3937
rect 336 139 432 3821
rect 996 3678 1028 3681
rect 996 3643 1028 3646
rect 993 3522 996 3554
rect 1028 3522 1031 3554
rect 996 3270 1028 3273
rect 996 3235 1028 3238
rect 993 3108 996 3140
rect 1028 3108 1031 3140
rect 996 2888 1028 2891
rect 996 2853 1028 2856
rect 993 2712 996 2744
rect 1028 2712 1031 2744
rect 996 2474 1028 2477
rect 996 2439 1028 2442
rect 993 2312 996 2344
rect 1028 2312 1031 2344
rect 996 2074 1028 2077
rect 996 2039 1028 2042
rect 993 1906 996 1938
rect 1028 1906 1031 1938
rect 996 1675 1028 1678
rect 996 1640 1028 1643
rect 993 1515 996 1547
rect 1028 1515 1031 1547
rect 996 1297 1028 1300
rect 996 1262 1028 1265
rect 993 1111 996 1143
rect 1028 1111 1031 1143
rect 996 870 1028 873
rect 996 835 1028 838
rect 993 708 996 740
rect 1028 708 1031 740
rect 996 492 1028 495
rect 996 457 1028 460
rect 993 313 996 345
rect 1028 313 1031 345
rect 368 110 400 113
rect 993 87 996 119
rect 1028 87 1031 119
rect 368 75 400 78
rect 1060 -49 1156 4287
rect 1251 4158 1347 4436
rect 1252 119 1348 3863
rect 1252 88 1272 119
rect 1304 88 1348 119
rect 1272 84 1304 87
rect 1060 -139 1063 -49
rect 1153 -139 1156 -49
rect 1060 -166 1156 -139
rect 870 -262 1575 -166
<< via1 >>
rect 80 3648 112 3680
rect 80 3520 112 3552
rect 80 3242 112 3274
rect 80 3123 112 3155
rect 80 2841 112 2873
rect 80 2731 112 2763
rect 80 2439 112 2471
rect 80 2307 112 2339
rect 80 2038 112 2070
rect 80 1927 112 1959
rect 80 1645 112 1677
rect 80 1515 112 1547
rect 80 1245 112 1277
rect 80 1097 112 1129
rect 80 844 112 876
rect 80 717 112 749
rect 80 444 112 476
rect 80 322 112 354
rect 80 78 112 110
rect 996 4030 1028 4062
rect 996 3905 1028 3937
rect 996 3646 1028 3678
rect 996 3522 1028 3554
rect 996 3238 1028 3270
rect 996 3108 1028 3140
rect 996 2856 1028 2888
rect 996 2712 1028 2744
rect 996 2442 1028 2474
rect 996 2312 1028 2344
rect 996 2042 1028 2074
rect 996 1906 1028 1938
rect 996 1643 1028 1675
rect 996 1515 1028 1547
rect 996 1265 1028 1297
rect 996 1111 1028 1143
rect 996 838 1028 870
rect 996 708 1028 740
rect 996 460 1028 492
rect 996 313 1028 345
rect 368 78 400 110
rect 996 87 1028 119
rect 1272 87 1304 119
<< metal2 >>
rect 993 4030 996 4062
rect 1028 4030 1031 4062
rect 996 3937 1028 4030
rect 996 3902 1028 3905
rect 77 3648 80 3680
rect 112 3648 115 3680
rect 80 3552 112 3648
rect 993 3646 996 3678
rect 1028 3646 1031 3678
rect 80 3517 112 3520
rect 996 3554 1028 3646
rect 996 3519 1028 3522
rect 77 3242 80 3274
rect 112 3242 115 3274
rect 80 3155 112 3242
rect 993 3238 996 3270
rect 1028 3238 1031 3270
rect 80 3120 112 3123
rect 996 3140 1028 3238
rect 996 3105 1028 3108
rect 77 2841 80 2873
rect 112 2841 115 2873
rect 993 2856 996 2888
rect 1028 2856 1031 2888
rect 80 2763 112 2841
rect 80 2728 112 2731
rect 996 2744 1028 2856
rect 996 2709 1028 2712
rect 77 2439 80 2471
rect 112 2439 115 2471
rect 993 2442 996 2474
rect 1028 2442 1031 2474
rect 80 2339 112 2439
rect 996 2344 1028 2442
rect 996 2309 1028 2312
rect 80 2304 112 2307
rect 77 2038 80 2070
rect 112 2038 115 2070
rect 993 2042 996 2074
rect 1028 2042 1031 2074
rect 80 1959 112 2038
rect 80 1924 112 1927
rect 996 1938 1028 2042
rect 996 1903 1028 1906
rect 77 1645 80 1677
rect 112 1645 115 1677
rect 80 1547 112 1645
rect 993 1643 996 1675
rect 1028 1643 1031 1675
rect 80 1512 112 1515
rect 996 1547 1028 1643
rect 996 1512 1028 1515
rect 77 1245 80 1277
rect 112 1245 115 1277
rect 993 1265 996 1297
rect 1028 1265 1031 1297
rect 80 1129 112 1245
rect 996 1143 1028 1265
rect 996 1108 1028 1111
rect 80 1094 112 1097
rect 77 844 80 876
rect 112 844 115 876
rect 80 749 112 844
rect 993 838 996 870
rect 1028 838 1031 870
rect 80 714 112 717
rect 996 740 1028 838
rect 996 705 1028 708
rect 77 444 80 476
rect 112 444 115 476
rect 993 460 996 492
rect 1028 460 1031 492
rect 80 354 112 444
rect 80 319 112 322
rect 996 345 1028 460
rect 996 310 1028 313
rect 996 119 1028 122
rect 80 110 112 113
rect 112 78 368 110
rect 400 78 403 110
rect 1028 87 1272 119
rect 1304 87 1307 119
rect 996 84 1028 87
rect 80 75 112 78
use JNWATR_PCH_4C5F0  xa2_0 ~/pro/aicex/ip/jnw_gr04_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 0 0 1 0
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_1
timestamp 1734044400
transform 1 0 0 0 1 400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_2
timestamp 1734044400
transform 1 0 0 0 1 800
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_3
timestamp 1734044400
transform 1 0 0 0 1 1200
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_4
timestamp 1734044400
transform 1 0 0 0 1 1600
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_5
timestamp 1734044400
transform 1 0 0 0 1 2000
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_6
timestamp 1734044400
transform 1 0 0 0 1 2400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_7
timestamp 1734044400
transform 1 0 0 0 1 2800
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_8
timestamp 1734044400
transform 1 0 0 0 1 3200
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2_9
timestamp 1734044400
transform 1 0 0 0 1 3600
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa3
timestamp 1734044400
transform 1 0 0 0 1 4000
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 916 0 1 0
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_1
timestamp 1734044400
transform 1 0 916 0 1 400
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_2
timestamp 1734044400
transform 1 0 916 0 1 800
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_3
timestamp 1734044400
transform 1 0 916 0 1 1200
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_4
timestamp 1734044400
transform 1 0 916 0 1 1600
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_5
timestamp 1734044400
transform 1 0 916 0 1 2000
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_6
timestamp 1734044400
transform 1 0 916 0 1 2400
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_7
timestamp 1734044400
transform 1 0 916 0 1 2800
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_8
timestamp 1734044400
transform 1 0 916 0 1 3200
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb1_9
timestamp 1734044400
transform 1 0 916 0 1 3600
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xb4
timestamp 1734044400
transform 1 0 916 0 1 4000
box -92 -64 668 464
<< labels >>
flabel metal1 157 4551 223 4637 0 FreeSans 800 0 0 0 VDD_1V8
port 1 nsew
flabel metal1 1088 -254 1154 -168 0 FreeSans 800 0 0 0 VSS
port 3 nsew
flabel metal1 1269 3495 1333 3722 0 FreeSans 800 0 0 0 I_IN
port 6 nsew
flabel metal1 354 4238 433 4296 0 FreeSans 800 0 0 0 I_OUT
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1492 4400
<< end >>
