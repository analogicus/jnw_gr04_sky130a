magic
tech sky130A
magscale 1 2
timestamp 1744566163
<< locali >>
rect -96 8882 298 9074
rect 478 8882 1242 9074
rect -96 8618 96 8882
rect 1050 8714 1242 8882
rect 1736 -102 1928 164
rect 1736 -278 2126 -102
rect 2882 -102 3074 76
rect 2306 -278 3074 -102
rect 1736 -294 3074 -278
<< viali >>
rect 298 8882 478 9074
rect 2126 -278 2306 -98
<< metal1 >>
rect -204 9126 1274 9318
rect 288 9086 480 9126
rect 288 9074 484 9086
rect 288 8882 298 9074
rect 478 8882 484 9074
rect 288 8870 484 8882
rect 1412 8872 2694 9064
rect 160 8168 224 8174
rect 160 7882 224 8135
rect 160 7360 224 7366
rect 160 7290 224 7296
rect 154 7040 160 7104
rect 224 7040 230 7104
rect 160 6548 224 6554
rect 160 6478 224 6484
rect 154 6246 160 6310
rect 224 6246 230 6310
rect 160 5746 224 5752
rect 160 5676 224 5682
rect 154 5462 160 5526
rect 224 5462 230 5526
rect 160 4942 224 4948
rect 160 4872 224 4878
rect 154 4614 160 4678
rect 224 4614 230 4678
rect 160 4140 224 4146
rect 160 4070 224 4076
rect 154 3854 160 3918
rect 224 3854 230 3918
rect 160 3354 224 3360
rect 160 3284 224 3290
rect 154 3030 160 3094
rect 224 3030 230 3094
rect 160 2554 224 2560
rect 160 2484 224 2490
rect 154 2194 160 2258
rect 224 2194 230 2258
rect 160 1752 224 1758
rect 160 1682 224 1688
rect 154 1434 160 1498
rect 224 1434 230 1498
rect 160 952 224 958
rect 160 882 224 888
rect 154 644 160 708
rect 224 644 230 708
rect 154 156 160 220
rect 224 156 230 220
rect 288 24 480 8870
rect 672 8438 976 8630
rect 1412 7834 1604 8872
rect 1992 8124 2056 8130
rect 1992 8054 2056 8060
rect 672 7642 1638 7834
rect 1986 7810 1992 7874
rect 2056 7810 2062 7874
rect 672 278 864 7642
rect 1992 7356 2056 7362
rect 1992 7286 2056 7292
rect 1986 7044 1992 7108
rect 2056 7044 2062 7108
rect 1992 6540 2056 6546
rect 1992 6470 2056 6476
rect 1986 6216 1992 6280
rect 2056 6216 2062 6280
rect 1992 5776 2056 5782
rect 1992 5706 2056 5712
rect 1986 5424 1992 5488
rect 2056 5424 2062 5488
rect 1992 4948 2056 4954
rect 1992 4878 2056 4884
rect 1986 4624 1992 4688
rect 2056 4624 2062 4688
rect 1992 4148 2056 4154
rect 1992 4078 2056 4084
rect 1986 3812 1992 3876
rect 2056 3812 2062 3876
rect 1992 3350 2056 3356
rect 1992 3280 2056 3286
rect 1986 3030 1992 3094
rect 2056 3030 2062 3094
rect 1992 2594 2056 2600
rect 1992 2524 2056 2530
rect 1986 2222 1992 2286
rect 2056 2222 2062 2286
rect 1992 1740 2056 1746
rect 1992 1670 2056 1676
rect 1986 1416 1992 1480
rect 2056 1416 2062 1480
rect 1992 984 2056 990
rect 1992 914 2056 920
rect 1986 626 1992 690
rect 2056 626 2062 690
rect 736 220 800 226
rect 1986 174 1992 238
rect 2056 174 2062 238
rect 736 150 800 156
rect 2120 -98 2312 8574
rect 2502 8316 2694 8872
rect 2504 238 2696 7726
rect 2504 176 2544 238
rect 2608 176 2696 238
rect 2544 168 2608 174
rect 2120 -278 2126 -98
rect 2306 -278 2312 -98
rect 2120 -332 2312 -278
rect 1740 -524 3150 -332
<< via1 >>
rect 160 7296 224 7360
rect 160 7040 224 7104
rect 160 6484 224 6548
rect 160 6246 224 6310
rect 160 5682 224 5746
rect 160 5462 224 5526
rect 160 4878 224 4942
rect 160 4614 224 4678
rect 160 4076 224 4140
rect 160 3854 224 3918
rect 160 3290 224 3354
rect 160 3030 224 3094
rect 160 2490 224 2554
rect 160 2194 224 2258
rect 160 1688 224 1752
rect 160 1434 224 1498
rect 160 888 224 952
rect 160 644 224 708
rect 160 156 224 220
rect 1992 8060 2056 8124
rect 1992 7810 2056 7874
rect 1992 7292 2056 7356
rect 1992 7044 2056 7108
rect 1992 6476 2056 6540
rect 1992 6216 2056 6280
rect 1992 5712 2056 5776
rect 1992 5424 2056 5488
rect 1992 4884 2056 4948
rect 1992 4624 2056 4688
rect 1992 4084 2056 4148
rect 1992 3812 2056 3876
rect 1992 3286 2056 3350
rect 1992 3030 2056 3094
rect 1992 2530 2056 2594
rect 1992 2222 2056 2286
rect 1992 1676 2056 1740
rect 1992 1416 2056 1480
rect 1992 920 2056 984
rect 1992 626 2056 690
rect 736 156 800 220
rect 1992 174 2056 238
rect 2544 174 2608 238
<< metal2 >>
rect 1986 8060 1992 8124
rect 2056 8060 2062 8124
rect 1992 7874 2056 8060
rect 1992 7804 2056 7810
rect 154 7296 160 7360
rect 224 7296 230 7360
rect 160 7104 224 7296
rect 1986 7292 1992 7356
rect 2056 7292 2062 7356
rect 160 7034 224 7040
rect 1992 7108 2056 7292
rect 1992 7038 2056 7044
rect 154 6484 160 6548
rect 224 6484 230 6548
rect 160 6310 224 6484
rect 1986 6476 1992 6540
rect 2056 6476 2062 6540
rect 160 6240 224 6246
rect 1992 6280 2056 6476
rect 1992 6210 2056 6216
rect 154 5682 160 5746
rect 224 5682 230 5746
rect 1986 5712 1992 5776
rect 2056 5712 2062 5776
rect 160 5526 224 5682
rect 160 5456 224 5462
rect 1992 5488 2056 5712
rect 1992 5418 2056 5424
rect 154 4878 160 4942
rect 224 4878 230 4942
rect 1986 4884 1992 4948
rect 2056 4884 2062 4948
rect 160 4678 224 4878
rect 1992 4688 2056 4884
rect 1992 4618 2056 4624
rect 160 4608 224 4614
rect 154 4076 160 4140
rect 224 4076 230 4140
rect 1986 4084 1992 4148
rect 2056 4084 2062 4148
rect 160 3918 224 4076
rect 160 3848 224 3854
rect 1992 3876 2056 4084
rect 1992 3806 2056 3812
rect 154 3290 160 3354
rect 224 3290 230 3354
rect 160 3094 224 3290
rect 1986 3286 1992 3350
rect 2056 3286 2062 3350
rect 160 3024 224 3030
rect 1992 3094 2056 3286
rect 1992 3024 2056 3030
rect 154 2490 160 2554
rect 224 2490 230 2554
rect 1986 2530 1992 2594
rect 2056 2530 2062 2594
rect 160 2258 224 2490
rect 1992 2286 2056 2530
rect 1992 2216 2056 2222
rect 160 2188 224 2194
rect 154 1688 160 1752
rect 224 1688 230 1752
rect 160 1498 224 1688
rect 1986 1676 1992 1740
rect 2056 1676 2062 1740
rect 160 1428 224 1434
rect 1992 1480 2056 1676
rect 1992 1410 2056 1416
rect 154 888 160 952
rect 224 888 230 952
rect 1986 920 1992 984
rect 2056 920 2062 984
rect 160 708 224 888
rect 160 638 224 644
rect 1992 690 2056 920
rect 1992 620 2056 626
rect 1992 238 2056 244
rect 160 220 224 226
rect 224 156 736 220
rect 800 156 806 220
rect 2056 174 2544 238
rect 2608 174 2614 238
rect 1992 168 2056 174
rect 160 150 224 156
use JNWATR_PCH_4C5F0__0  xa2_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_1
timestamp 1734044400
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_2
timestamp 1734044400
transform 1 0 0 0 1 1600
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_3
timestamp 1734044400
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_4
timestamp 1734044400
transform 1 0 0 0 1 3200
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_5
timestamp 1734044400
transform 1 0 0 0 1 4000
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_6
timestamp 1734044400
transform 1 0 0 0 1 4800
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_7
timestamp 1734044400
transform 1 0 0 0 1 5600
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_8
timestamp 1734044400
transform 1 0 0 0 1 6400
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa2_9
timestamp 1734044400
transform 1 0 0 0 1 7200
box -184 -128 1336 928
use JNWATR_PCH_4C5F0__0  xa3
timestamp 1734044400
transform 1 0 0 0 1 8000
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 1832 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_1
timestamp 1734044400
transform 1 0 1832 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_2
timestamp 1734044400
transform 1 0 1832 0 1 1600
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_3
timestamp 1734044400
transform 1 0 1832 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_4
timestamp 1734044400
transform 1 0 1832 0 1 3200
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_5
timestamp 1734044400
transform 1 0 1832 0 1 4000
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_6
timestamp 1734044400
transform 1 0 1832 0 1 4800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_7
timestamp 1734044400
transform 1 0 1832 0 1 5600
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_8
timestamp 1734044400
transform 1 0 1832 0 1 6400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb1_9
timestamp 1734044400
transform 1 0 1832 0 1 7200
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xb4
timestamp 1734044400
transform 1 0 1832 0 1 8000
box -184 -128 1336 928
<< labels >>
flabel metal1 314 9102 446 9274 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel metal1 2176 -508 2308 -336 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal1 2538 6990 2666 7444 0 FreeSans 1600 0 0 0 I_IN
port 6 nsew
flabel metal1 708 8476 866 8592 0 FreeSans 1600 0 0 0 I_OUT
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 2984 8800
<< end >>
