*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/Opamp_lpe.spi
#else
.include ../../../work/xsch/Opamp.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param AVDD = {vdda}
.param VCM = {AVDD * 0.5}  
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  VSS  dc {AVDD}
VSS  VSS  0    dc 0

* Biasing the non-inverting input to a DC common-mode voltage
Vcm VIP VSS  dc {VCM}

* Small-signal AC source at inverting input
Vac  VIN  VSS  ac 1mV

*-----------------------------------------------------------------
* DUT (Open-loop configuration)
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
*.save v(Vo) v(VIP) v(VIN)
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit 

tran 10n 10u


* AC Analysis: Sweep frequency from 1 Hz to 1 GHz
*ac dec 100 1 1G
*plot v(Vo) v(VIN)

write 

quit
.endc

.end
