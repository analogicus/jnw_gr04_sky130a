*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR04_lpe.spi
#else
.include ../../../work/xsch/JNW_GR04.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}
.param PERIOD_CLK = 48n
.param PW_CLK = PERIOD_CLK/2


*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VCLK clk 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names
VB0 b.0 b<0> dc 0
VB1 b.1 b<1> dc 0
VB2 b.2 b<2> dc 0
VB3 b.3 b<3> dc 0
VB4 b.4 b<4> dc 0
VB5 b.5 b<5> dc 0
VB6 b.6 b<6> dc 0
VB7 b.7 b<7> dc 0

VOUT analog_out OUT dc 0

*-----------------------------------------------------------------
* Testbench for comparator functionality
*-----------------------------------------------------------------
* Generate a pulse signal on INP to test the comparator's behavior
*Vin INP 0 DC 0V PULSE (0V 1.8V 0 10n 10n 50n 100n)  
* Generate a pulse from 0V to 1.8V with a longer high time

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit



*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )




set fend = .raw
*foreach vtemp -40 -35 -30 -25 -20 -15 -10 -5 0 5 10 15 20 25 30 35 40 45 50 55 60 65 70 75 80 85 90 95 100 105 110 115 120
*foreach vtemp -40 -20 0 20 40 60 80 100 120
foreach vtemp -40 0 40 80 120
*foreach vtemp 80
  option temp=$vtemp
  tran 1n 30u 1p
  write {cicname}_$vtemp$fend
end

* Output results
*write
quit

.endc

.end
