magic
tech sky130A
magscale 1 2
timestamp 1744383272
<< viali >>
rect 7021 8925 7055 8959
rect 7941 8925 7975 8959
rect 7205 8789 7239 8823
rect 7389 8789 7423 8823
rect 4629 8517 4663 8551
rect 4845 8517 4879 8551
rect 1685 8449 1719 8483
rect 2053 8449 2087 8483
rect 4537 8449 4571 8483
rect 6101 8449 6135 8483
rect 3157 8381 3191 8415
rect 4261 8381 4295 8415
rect 4445 8381 4479 8415
rect 7205 8381 7239 8415
rect 7941 8381 7975 8415
rect 1501 8313 1535 8347
rect 1869 8313 1903 8347
rect 4353 8313 4387 8347
rect 4997 8313 5031 8347
rect 7389 8313 7423 8347
rect 2605 8245 2639 8279
rect 4813 8245 4847 8279
rect 6653 8245 6687 8279
rect 2421 8041 2455 8075
rect 4997 8041 5031 8075
rect 7757 8041 7791 8075
rect 3065 7905 3099 7939
rect 5181 7905 5215 7939
rect 5733 7905 5767 7939
rect 6377 7905 6411 7939
rect 1685 7837 1719 7871
rect 3985 7837 4019 7871
rect 4537 7837 4571 7871
rect 5273 7837 5307 7871
rect 5365 7837 5399 7871
rect 5457 7837 5491 7871
rect 6644 7837 6678 7871
rect 2329 7769 2363 7803
rect 2881 7769 2915 7803
rect 2789 7701 2823 7735
rect 6285 7701 6319 7735
rect 1501 7497 1535 7531
rect 7757 7497 7791 7531
rect 2614 7429 2648 7463
rect 3218 7429 3252 7463
rect 6101 7429 6135 7463
rect 6644 7429 6678 7463
rect 4445 7361 4479 7395
rect 6377 7361 6411 7395
rect 2881 7293 2915 7327
rect 2973 7293 3007 7327
rect 4353 7157 4387 7191
rect 6193 6953 6227 6987
rect 2973 6817 3007 6851
rect 4353 6817 4387 6851
rect 7113 6817 7147 6851
rect 7205 6817 7239 6851
rect 3341 6749 3375 6783
rect 3617 6749 3651 6783
rect 4813 6749 4847 6783
rect 6561 6749 6595 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 2728 6681 2762 6715
rect 3525 6681 3559 6715
rect 4169 6681 4203 6715
rect 5080 6681 5114 6715
rect 7573 6681 7607 6715
rect 1593 6613 1627 6647
rect 3157 6613 3191 6647
rect 3801 6613 3835 6647
rect 4261 6613 4295 6647
rect 6377 6613 6411 6647
rect 6653 6613 6687 6647
rect 7021 6613 7055 6647
rect 2789 6409 2823 6443
rect 5917 6409 5951 6443
rect 6009 6409 6043 6443
rect 6193 6409 6227 6443
rect 7021 6409 7055 6443
rect 7481 6409 7515 6443
rect 7113 6341 7147 6375
rect 2145 6273 2179 6307
rect 2881 6273 2915 6307
rect 3148 6273 3182 6307
rect 4445 6273 4479 6307
rect 4537 6273 4571 6307
rect 4997 6273 5031 6307
rect 5153 6273 5187 6307
rect 5411 6273 5445 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 7757 6273 7791 6307
rect 4813 6205 4847 6239
rect 5267 6205 5301 6239
rect 6193 6205 6227 6239
rect 6837 6205 6871 6239
rect 7941 6205 7975 6239
rect 4721 6137 4755 6171
rect 6377 6137 6411 6171
rect 4261 6069 4295 6103
rect 4905 6069 4939 6103
rect 5733 6069 5767 6103
rect 7573 6069 7607 6103
rect 2697 5865 2731 5899
rect 2973 5865 3007 5899
rect 3893 5865 3927 5899
rect 7297 5865 7331 5899
rect 2421 5797 2455 5831
rect 2881 5797 2915 5831
rect 3617 5729 3651 5763
rect 7389 5729 7423 5763
rect 2145 5661 2179 5695
rect 2237 5661 2271 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 5917 5661 5951 5695
rect 8033 5661 8067 5695
rect 2421 5593 2455 5627
rect 2513 5593 2547 5627
rect 6162 5593 6196 5627
rect 2723 5525 2757 5559
rect 5365 5525 5399 5559
rect 2513 5321 2547 5355
rect 6377 5321 6411 5355
rect 2145 5253 2179 5287
rect 2361 5253 2395 5287
rect 2973 5253 3007 5287
rect 7941 5253 7975 5287
rect 1777 5185 1811 5219
rect 2789 5185 2823 5219
rect 3065 5185 3099 5219
rect 3617 5185 3651 5219
rect 4721 5185 4755 5219
rect 5549 5185 5583 5219
rect 7021 5185 7055 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 3249 5117 3283 5151
rect 3341 5117 3375 5151
rect 3801 5117 3835 5151
rect 4445 5117 4479 5151
rect 4905 5117 4939 5151
rect 7665 5117 7699 5151
rect 1961 5049 1995 5083
rect 5457 5049 5491 5083
rect 2329 4981 2363 5015
rect 2605 4981 2639 5015
rect 4629 4981 4663 5015
rect 6193 4981 6227 5015
rect 7113 4981 7147 5015
rect 1961 4777 1995 4811
rect 3801 4777 3835 4811
rect 6837 4777 6871 4811
rect 1685 4709 1719 4743
rect 2973 4641 3007 4675
rect 7389 4641 7423 4675
rect 1409 4573 1443 4607
rect 2237 4573 2271 4607
rect 3525 4573 3559 4607
rect 4353 4573 4387 4607
rect 4721 4573 4755 4607
rect 5365 4573 5399 4607
rect 7757 4573 7791 4607
rect 1685 4505 1719 4539
rect 1777 4505 1811 4539
rect 1993 4505 2027 4539
rect 5632 4505 5666 4539
rect 7297 4505 7331 4539
rect 1501 4437 1535 4471
rect 2145 4437 2179 4471
rect 2881 4437 2915 4471
rect 5273 4437 5307 4471
rect 6745 4437 6779 4471
rect 7205 4437 7239 4471
rect 7941 4437 7975 4471
rect 6101 4233 6135 4267
rect 7757 4233 7791 4267
rect 2666 4165 2700 4199
rect 5006 4097 5040 4131
rect 5457 4097 5491 4131
rect 6644 4097 6678 4131
rect 1777 4029 1811 4063
rect 2421 4029 2455 4063
rect 5273 4029 5307 4063
rect 6377 4029 6411 4063
rect 3801 3961 3835 3995
rect 2329 3893 2363 3927
rect 3893 3893 3927 3927
rect 1593 3689 1627 3723
rect 3341 3621 3375 3655
rect 3893 3621 3927 3655
rect 5641 3621 5675 3655
rect 7849 3621 7883 3655
rect 1961 3553 1995 3587
rect 1593 3485 1627 3519
rect 1869 3485 1903 3519
rect 4261 3485 4295 3519
rect 4353 3485 4387 3519
rect 6193 3485 6227 3519
rect 6449 3485 6483 3519
rect 7665 3485 7699 3519
rect 2206 3417 2240 3451
rect 1777 3349 1811 3383
rect 3801 3349 3835 3383
rect 7573 3349 7607 3383
rect 1593 3145 1627 3179
rect 3525 3145 3559 3179
rect 3985 3145 4019 3179
rect 4537 3145 4571 3179
rect 7757 3145 7791 3179
rect 2706 3009 2740 3043
rect 2973 3009 3007 3043
rect 3249 3009 3283 3043
rect 3617 3009 3651 3043
rect 3709 3009 3743 3043
rect 4169 3009 4203 3043
rect 5650 3009 5684 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 6193 3009 6227 3043
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 4077 2941 4111 2975
rect 4445 2941 4479 2975
rect 3341 2873 3375 2907
rect 3249 2805 3283 2839
rect 1685 2601 1719 2635
rect 2421 2601 2455 2635
rect 6193 2601 6227 2635
rect 6561 2601 6595 2635
rect 7573 2601 7607 2635
rect 3801 2533 3835 2567
rect 6745 2533 6779 2567
rect 7665 2533 7699 2567
rect 2329 2465 2363 2499
rect 2881 2465 2915 2499
rect 3065 2465 3099 2499
rect 4261 2465 4295 2499
rect 4445 2465 4479 2499
rect 5641 2465 5675 2499
rect 7205 2465 7239 2499
rect 7389 2465 7423 2499
rect 2789 2397 2823 2431
rect 3617 2397 3651 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 4905 2397 4939 2431
rect 6377 2397 6411 2431
rect 7113 2397 7147 2431
rect 8033 2397 8067 2431
rect 3433 2261 3467 2295
<< metal1 >>
rect 1104 9274 8372 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 8372 9274
rect 1104 9200 8372 9222
rect 7006 8916 7012 8968
rect 7064 8916 7070 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 7800 8928 7941 8956
rect 7800 8916 7806 8928
rect 7929 8925 7941 8928
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 7190 8780 7196 8832
rect 7248 8780 7254 8832
rect 7374 8780 7380 8832
rect 7432 8780 7438 8832
rect 1104 8730 8372 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8372 8730
rect 1104 8656 8372 8678
rect 4617 8551 4675 8557
rect 4617 8548 4629 8551
rect 4264 8520 4629 8548
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2130 8480 2136 8492
rect 2087 8452 2136 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 3142 8372 3148 8424
rect 3200 8372 3206 8424
rect 4264 8421 4292 8520
rect 4617 8517 4629 8520
rect 4663 8517 4675 8551
rect 4617 8511 4675 8517
rect 4833 8551 4891 8557
rect 4833 8517 4845 8551
rect 4879 8548 4891 8551
rect 6178 8548 6184 8560
rect 4879 8520 6184 8548
rect 4879 8517 4891 8520
rect 4833 8511 4891 8517
rect 6178 8508 6184 8520
rect 6236 8508 6242 8560
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4706 8480 4712 8492
rect 4571 8452 4712 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 6086 8440 6092 8492
rect 6144 8440 6150 8492
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 5350 8412 5356 8424
rect 4479 8384 5356 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 1854 8304 1860 8356
rect 1912 8304 1918 8356
rect 2590 8236 2596 8288
rect 2648 8236 2654 8288
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 4264 8276 4292 8375
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 6972 8384 7205 8412
rect 6972 8372 6978 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 7926 8372 7932 8424
rect 7984 8372 7990 8424
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 4614 8344 4620 8356
rect 4387 8316 4620 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 4985 8347 5043 8353
rect 4985 8313 4997 8347
rect 5031 8344 5043 8347
rect 5258 8344 5264 8356
rect 5031 8316 5264 8344
rect 5031 8313 5043 8316
rect 4985 8307 5043 8313
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 6730 8304 6736 8356
rect 6788 8344 6794 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 6788 8316 7389 8344
rect 6788 8304 6794 8316
rect 7377 8313 7389 8316
rect 7423 8313 7435 8347
rect 7377 8307 7435 8313
rect 3384 8248 4292 8276
rect 3384 8236 3390 8248
rect 4798 8236 4804 8288
rect 4856 8236 4862 8288
rect 6638 8236 6644 8288
rect 6696 8236 6702 8288
rect 1104 8186 8372 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 8372 8186
rect 1104 8112 8372 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 3142 8072 3148 8084
rect 2455 8044 3148 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 4856 8044 4997 8072
rect 4856 8032 4862 8044
rect 4985 8041 4997 8044
rect 5031 8041 5043 8075
rect 7006 8072 7012 8084
rect 4985 8035 5043 8041
rect 5736 8044 7012 8072
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3326 7936 3332 7948
rect 3099 7908 3332 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 4706 7936 4712 7948
rect 3988 7908 4712 7936
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 3988 7877 4016 7908
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5626 7936 5632 7948
rect 5215 7908 5632 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5736 7945 5764 8044
rect 7006 8032 7012 8044
rect 7064 8072 7070 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7064 8044 7757 8072
rect 7064 8032 7070 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 6144 7908 6377 7936
rect 6144 7896 6150 7908
rect 6365 7905 6377 7908
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 2280 7840 3985 7868
rect 2280 7828 2286 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 2317 7803 2375 7809
rect 2317 7769 2329 7803
rect 2363 7800 2375 7803
rect 2869 7803 2927 7809
rect 2869 7800 2881 7803
rect 2363 7772 2881 7800
rect 2363 7769 2375 7772
rect 2317 7763 2375 7769
rect 2869 7769 2881 7772
rect 2915 7769 2927 7803
rect 5276 7800 5304 7831
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5902 7868 5908 7880
rect 5491 7840 5908 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6638 7877 6644 7880
rect 6632 7868 6644 7877
rect 6599 7840 6644 7868
rect 6632 7831 6644 7840
rect 6638 7828 6644 7831
rect 6696 7828 6702 7880
rect 5276 7772 5488 7800
rect 2869 7763 2927 7769
rect 5460 7744 5488 7772
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 3234 7732 3240 7744
rect 2823 7704 3240 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 5442 7692 5448 7744
rect 5500 7692 5506 7744
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 7098 7732 7104 7744
rect 6319 7704 7104 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 1104 7642 8372 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8372 7642
rect 1104 7568 8372 7590
rect 1489 7531 1547 7537
rect 1489 7497 1501 7531
rect 1535 7528 1547 7531
rect 1670 7528 1676 7540
rect 1535 7500 1676 7528
rect 1535 7497 1547 7500
rect 1489 7491 1547 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 2590 7420 2596 7472
rect 2648 7469 2654 7472
rect 2648 7460 2660 7469
rect 2648 7432 2693 7460
rect 2648 7423 2660 7432
rect 2648 7420 2654 7423
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 3206 7463 3264 7469
rect 3206 7460 3218 7463
rect 2924 7432 3218 7460
rect 2924 7420 2930 7432
rect 3206 7429 3218 7432
rect 3252 7429 3264 7463
rect 3206 7423 3264 7429
rect 6086 7420 6092 7472
rect 6144 7420 6150 7472
rect 6632 7463 6690 7469
rect 6632 7429 6644 7463
rect 6678 7460 6690 7463
rect 6730 7460 6736 7472
rect 6678 7432 6736 7460
rect 6678 7429 6690 7432
rect 6632 7423 6690 7429
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 5350 7392 5356 7404
rect 4479 7364 5356 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 6104 7392 6132 7420
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6104 7364 6377 7392
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 2958 7324 2964 7336
rect 2915 7296 2964 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4522 7188 4528 7200
rect 4387 7160 4528 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4522 7148 4528 7160
rect 4580 7188 4586 7200
rect 4706 7188 4712 7200
rect 4580 7160 4712 7188
rect 4580 7148 4586 7160
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 1104 7098 8372 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 8372 7098
rect 1104 7024 8372 7046
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6181 6987 6239 6993
rect 6181 6984 6193 6987
rect 5960 6956 6193 6984
rect 5960 6944 5966 6956
rect 6181 6953 6193 6956
rect 6227 6953 6239 6987
rect 6181 6947 6239 6953
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 3384 6888 4384 6916
rect 3384 6876 3390 6888
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 4356 6857 4384 6888
rect 4341 6851 4399 6857
rect 3016 6820 3740 6848
rect 3016 6808 3022 6820
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 3292 6752 3341 6780
rect 3292 6740 3298 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3602 6740 3608 6792
rect 3660 6740 3666 6792
rect 3712 6780 3740 6820
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 6196 6848 6224 6947
rect 6822 6876 6828 6928
rect 6880 6916 6886 6928
rect 6880 6888 7236 6916
rect 6880 6876 6886 6888
rect 7006 6848 7012 6860
rect 6196 6820 7012 6848
rect 4341 6811 4399 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7098 6808 7104 6860
rect 7156 6808 7162 6860
rect 7208 6857 7236 6888
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6817 7251 6851
rect 7193 6811 7251 6817
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 3712 6752 4813 6780
rect 4801 6749 4813 6752
rect 4847 6780 4859 6783
rect 5994 6780 6000 6792
rect 4847 6752 6000 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 7650 6780 7656 6792
rect 6595 6752 7656 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 7834 6740 7840 6792
rect 7892 6740 7898 6792
rect 2716 6715 2774 6721
rect 2716 6681 2728 6715
rect 2762 6712 2774 6715
rect 3050 6712 3056 6724
rect 2762 6684 3056 6712
rect 2762 6681 2774 6684
rect 2716 6675 2774 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 3559 6684 4169 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 4157 6681 4169 6684
rect 4203 6712 4215 6715
rect 4706 6712 4712 6724
rect 4203 6684 4712 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 4706 6672 4712 6684
rect 4764 6712 4770 6724
rect 5068 6715 5126 6721
rect 4764 6684 4936 6712
rect 4764 6672 4770 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2130 6644 2136 6656
rect 1627 6616 2136 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 2648 6616 3157 6644
rect 2648 6604 2654 6616
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3145 6607 3203 6613
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3660 6616 3801 6644
rect 3660 6604 3666 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4246 6604 4252 6656
rect 4304 6604 4310 6656
rect 4908 6644 4936 6684
rect 5068 6681 5080 6715
rect 5114 6712 5126 6715
rect 5258 6712 5264 6724
rect 5114 6684 5264 6712
rect 5114 6681 5126 6684
rect 5068 6675 5126 6681
rect 5258 6672 5264 6684
rect 5316 6672 5322 6724
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 7561 6715 7619 6721
rect 7561 6712 7573 6715
rect 5684 6684 7573 6712
rect 5684 6672 5690 6684
rect 7561 6681 7573 6684
rect 7607 6681 7619 6715
rect 7561 6675 7619 6681
rect 6270 6644 6276 6656
rect 4908 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6362 6604 6368 6656
rect 6420 6604 6426 6656
rect 6641 6647 6699 6653
rect 6641 6613 6653 6647
rect 6687 6644 6699 6647
rect 6914 6644 6920 6656
rect 6687 6616 6920 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7006 6604 7012 6656
rect 7064 6604 7070 6656
rect 1104 6554 8372 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8372 6554
rect 1104 6480 8372 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 4246 6440 4252 6452
rect 2823 6412 4252 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5074 6400 5080 6452
rect 5132 6400 5138 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5442 6440 5448 6452
rect 5224 6412 5448 6440
rect 5224 6400 5230 6412
rect 5442 6400 5448 6412
rect 5500 6440 5506 6452
rect 5902 6440 5908 6452
rect 5500 6412 5908 6440
rect 5500 6400 5506 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6086 6440 6092 6452
rect 6043 6412 6092 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6178 6400 6184 6452
rect 6236 6400 6242 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 7009 6443 7067 6449
rect 6328 6412 6960 6440
rect 6328 6400 6334 6412
rect 2406 6332 2412 6384
rect 2464 6372 2470 6384
rect 4614 6372 4620 6384
rect 2464 6344 4620 6372
rect 2464 6332 2470 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 2130 6264 2136 6316
rect 2188 6264 2194 6316
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 2958 6304 2964 6316
rect 2915 6276 2964 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3142 6313 3148 6316
rect 3136 6267 3148 6313
rect 3142 6264 3148 6267
rect 3200 6264 3206 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 4448 6236 4476 6267
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 4706 6264 4712 6316
rect 4764 6264 4770 6316
rect 4982 6264 4988 6316
rect 5040 6264 5046 6316
rect 5083 6304 5111 6400
rect 6454 6372 6460 6384
rect 5552 6344 6460 6372
rect 5442 6313 5448 6316
rect 5141 6307 5199 6313
rect 5141 6304 5153 6307
rect 5083 6276 5153 6304
rect 5141 6273 5153 6276
rect 5187 6273 5199 6307
rect 5141 6267 5199 6273
rect 5399 6307 5448 6313
rect 5399 6273 5411 6307
rect 5445 6273 5448 6307
rect 5399 6267 5448 6273
rect 5442 6264 5448 6267
rect 5500 6264 5506 6316
rect 5552 6313 5580 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5684 6276 5825 6304
rect 5684 6264 5690 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 6638 6264 6644 6316
rect 6696 6264 6702 6316
rect 6932 6304 6960 6412
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 7374 6440 7380 6452
rect 7055 6412 7380 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 7926 6440 7932 6452
rect 7515 6412 7932 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 7101 6375 7159 6381
rect 7101 6341 7113 6375
rect 7147 6372 7159 6375
rect 7834 6372 7840 6384
rect 7147 6344 7840 6372
rect 7147 6341 7159 6344
rect 7101 6335 7159 6341
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 6932 6276 7757 6304
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 4724 6236 4752 6264
rect 4448 6208 4752 6236
rect 4798 6196 4804 6248
rect 4856 6196 4862 6248
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 5255 6239 5313 6245
rect 5255 6236 5267 6239
rect 4948 6208 5267 6236
rect 4948 6196 4954 6208
rect 5255 6205 5267 6208
rect 5301 6205 5313 6239
rect 5255 6199 5313 6205
rect 6178 6196 6184 6248
rect 6236 6196 6242 6248
rect 6822 6196 6828 6248
rect 6880 6196 6886 6248
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7156 6208 7941 6236
rect 7156 6196 7162 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 4709 6171 4767 6177
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 6365 6171 6423 6177
rect 6365 6168 6377 6171
rect 4755 6140 6377 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 6365 6137 6377 6140
rect 6411 6137 6423 6171
rect 6365 6131 6423 6137
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3970 6100 3976 6112
rect 3292 6072 3976 6100
rect 3292 6060 3298 6072
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 4028 6072 4261 6100
rect 4028 6060 4034 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4893 6103 4951 6109
rect 4893 6069 4905 6103
rect 4939 6100 4951 6103
rect 5258 6100 5264 6112
rect 4939 6072 5264 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5718 6060 5724 6112
rect 5776 6060 5782 6112
rect 5902 6060 5908 6112
rect 5960 6100 5966 6112
rect 6638 6100 6644 6112
rect 5960 6072 6644 6100
rect 5960 6060 5966 6072
rect 6638 6060 6644 6072
rect 6696 6100 6702 6112
rect 7561 6103 7619 6109
rect 7561 6100 7573 6103
rect 6696 6072 7573 6100
rect 6696 6060 6702 6072
rect 7561 6069 7573 6072
rect 7607 6069 7619 6103
rect 7561 6063 7619 6069
rect 1104 6010 8372 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 8372 6010
rect 1104 5936 8372 5958
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2648 5868 2697 5896
rect 2648 5856 2654 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 2958 5856 2964 5908
rect 3016 5856 3022 5908
rect 3142 5896 3148 5908
rect 3068 5868 3148 5896
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5828 2467 5831
rect 2774 5828 2780 5840
rect 2455 5800 2780 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 2869 5831 2927 5837
rect 2869 5797 2881 5831
rect 2915 5828 2927 5831
rect 3068 5828 3096 5868
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 4890 5896 4896 5908
rect 3936 5868 4896 5896
rect 3936 5856 3942 5868
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 7098 5896 7104 5908
rect 5000 5868 7104 5896
rect 2915 5800 3096 5828
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 3568 5800 3740 5828
rect 3568 5788 3574 5800
rect 2314 5760 2320 5772
rect 2148 5732 2320 5760
rect 2148 5701 2176 5732
rect 2314 5720 2320 5732
rect 2372 5760 2378 5772
rect 3528 5760 3556 5788
rect 2372 5732 3556 5760
rect 2372 5720 2378 5732
rect 3602 5720 3608 5772
rect 3660 5720 3666 5772
rect 3712 5760 3740 5800
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 5000 5828 5028 5868
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 7834 5896 7840 5908
rect 7331 5868 7840 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 4028 5800 5028 5828
rect 4028 5788 4034 5800
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 5902 5828 5908 5840
rect 5132 5800 5908 5828
rect 5132 5788 5138 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 7392 5769 7420 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 7377 5763 7435 5769
rect 3712 5732 4016 5760
rect 3988 5704 4016 5732
rect 7377 5729 7389 5763
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2222 5652 2228 5704
rect 2280 5652 2286 5704
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 2406 5584 2412 5636
rect 2464 5584 2470 5636
rect 2498 5584 2504 5636
rect 2556 5584 2562 5636
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 3804 5624 3832 5655
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 5994 5692 6000 5704
rect 5951 5664 6000 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6454 5652 6460 5704
rect 6512 5692 6518 5704
rect 8018 5692 8024 5704
rect 6512 5664 8024 5692
rect 6512 5652 6518 5664
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 5166 5624 5172 5636
rect 2924 5596 5172 5624
rect 2924 5584 2930 5596
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 5718 5584 5724 5636
rect 5776 5624 5782 5636
rect 6150 5627 6208 5633
rect 6150 5624 6162 5627
rect 5776 5596 6162 5624
rect 5776 5584 5782 5596
rect 6150 5593 6162 5596
rect 6196 5593 6208 5627
rect 6150 5587 6208 5593
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 7650 5624 7656 5636
rect 6420 5596 7656 5624
rect 6420 5584 6426 5596
rect 7650 5584 7656 5596
rect 7708 5584 7714 5636
rect 2711 5559 2769 5565
rect 2711 5525 2723 5559
rect 2757 5556 2769 5559
rect 3878 5556 3884 5568
rect 2757 5528 3884 5556
rect 2757 5525 2769 5528
rect 2711 5519 2769 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 5350 5516 5356 5568
rect 5408 5516 5414 5568
rect 1104 5466 8372 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8372 5466
rect 1104 5392 8372 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 4798 5352 4804 5364
rect 2547 5324 4804 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6236 5324 6377 5352
rect 6236 5312 6242 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 2038 5244 2044 5296
rect 2096 5284 2102 5296
rect 2133 5287 2191 5293
rect 2133 5284 2145 5287
rect 2096 5256 2145 5284
rect 2096 5244 2102 5256
rect 2133 5253 2145 5256
rect 2179 5253 2191 5287
rect 2133 5247 2191 5253
rect 2349 5287 2407 5293
rect 2349 5253 2361 5287
rect 2395 5284 2407 5287
rect 2866 5284 2872 5296
rect 2395 5256 2872 5284
rect 2395 5253 2407 5256
rect 2349 5247 2407 5253
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3510 5284 3516 5296
rect 3007 5256 3516 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 3896 5256 5580 5284
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2222 5216 2228 5228
rect 1811 5188 2228 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2774 5176 2780 5228
rect 2832 5176 2838 5228
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3896 5216 3924 5256
rect 3651 5188 3924 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 3068 5148 3096 5179
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4028 5188 4721 5216
rect 4028 5176 4034 5188
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 1728 5120 3096 5148
rect 1728 5108 1734 5120
rect 3234 5108 3240 5160
rect 3292 5108 3298 5160
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 2682 5080 2688 5092
rect 1995 5052 2688 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 2682 5040 2688 5052
rect 2740 5040 2746 5092
rect 3344 5080 3372 5111
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3476 5120 3801 5148
rect 3476 5108 3482 5120
rect 3789 5117 3801 5120
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4614 5148 4620 5160
rect 4479 5120 4620 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 3602 5080 3608 5092
rect 3344 5052 3608 5080
rect 3602 5040 3608 5052
rect 3660 5080 3666 5092
rect 4522 5080 4528 5092
rect 3660 5052 4528 5080
rect 3660 5040 3666 5052
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 3752 4984 4629 5012
rect 3752 4972 3758 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4617 4975 4675 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4816 5012 4844 5256
rect 5552 5225 5580 5256
rect 5902 5244 5908 5296
rect 5960 5284 5966 5296
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 5960 5256 7941 5284
rect 5960 5244 5966 5256
rect 7929 5253 7941 5256
rect 7975 5253 7987 5287
rect 7929 5247 7987 5253
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7834 5176 7840 5228
rect 7892 5176 7898 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5148 4951 5151
rect 6362 5148 6368 5160
rect 4939 5120 6368 5148
rect 4939 5117 4951 5120
rect 4893 5111 4951 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 5445 5083 5503 5089
rect 5445 5049 5457 5083
rect 5491 5080 5503 5083
rect 7190 5080 7196 5092
rect 5491 5052 7196 5080
rect 5491 5049 5503 5052
rect 5445 5043 5503 5049
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 4764 4984 4844 5012
rect 4764 4972 4770 4984
rect 6178 4972 6184 5024
rect 6236 4972 6242 5024
rect 6638 4972 6644 5024
rect 6696 5012 6702 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6696 4984 7113 5012
rect 6696 4972 6702 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 1104 4922 8372 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 8372 4922
rect 1104 4848 8372 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2590 4808 2596 4820
rect 1995 4780 2596 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2832 4780 3801 4808
rect 2832 4768 2838 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 6825 4811 6883 4817
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 7650 4808 7656 4820
rect 6871 4780 7656 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 1578 4700 1584 4752
rect 1636 4740 1642 4752
rect 1673 4743 1731 4749
rect 1673 4740 1685 4743
rect 1636 4712 1685 4740
rect 1636 4700 1642 4712
rect 1673 4709 1685 4712
rect 1719 4709 1731 4743
rect 2498 4740 2504 4752
rect 1673 4703 1731 4709
rect 1780 4712 2504 4740
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 1780 4604 1808 4712
rect 2498 4700 2504 4712
rect 2556 4740 2562 4752
rect 3050 4740 3056 4752
rect 2556 4712 3056 4740
rect 2556 4700 2562 4712
rect 3050 4700 3056 4712
rect 3108 4740 3114 4752
rect 3326 4740 3332 4752
rect 3108 4712 3332 4740
rect 3108 4700 3114 4712
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2056 4644 2973 4672
rect 2056 4604 2084 4644
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6880 4644 7389 4672
rect 6880 4632 6886 4644
rect 7377 4641 7389 4644
rect 7423 4672 7435 4675
rect 7650 4672 7656 4684
rect 7423 4644 7656 4672
rect 7423 4641 7435 4644
rect 7377 4635 7435 4641
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 1397 4567 1455 4573
rect 1596 4576 1808 4604
rect 1412 4536 1440 4567
rect 1596 4536 1624 4576
rect 1412 4508 1624 4536
rect 1670 4496 1676 4548
rect 1728 4496 1734 4548
rect 1780 4545 1808 4576
rect 1872 4576 2084 4604
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4505 1823 4539
rect 1765 4499 1823 4505
rect 1872 4480 1900 4576
rect 2222 4564 2228 4616
rect 2280 4564 2286 4616
rect 3510 4564 3516 4616
rect 3568 4564 3574 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4212 4576 4353 4604
rect 4212 4564 4218 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5442 4604 5448 4616
rect 5399 4576 5448 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 1981 4539 2039 4545
rect 1981 4505 1993 4539
rect 2027 4536 2039 4539
rect 3694 4536 3700 4548
rect 2027 4508 3700 4536
rect 2027 4505 2039 4508
rect 1981 4499 2039 4505
rect 3694 4496 3700 4508
rect 3752 4496 3758 4548
rect 4724 4536 4752 4567
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 7742 4604 7748 4616
rect 5552 4576 7748 4604
rect 5552 4536 5580 4576
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 4724 4508 5580 4536
rect 5620 4539 5678 4545
rect 5620 4505 5632 4539
rect 5666 4536 5678 4539
rect 6086 4536 6092 4548
rect 5666 4508 6092 4536
rect 5666 4505 5678 4508
rect 5620 4499 5678 4505
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 7285 4539 7343 4545
rect 7285 4536 7297 4539
rect 6288 4508 7297 4536
rect 1489 4471 1547 4477
rect 1489 4437 1501 4471
rect 1535 4468 1547 4471
rect 1854 4468 1860 4480
rect 1535 4440 1860 4468
rect 1535 4437 1547 4440
rect 1489 4431 1547 4437
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 2130 4428 2136 4480
rect 2188 4428 2194 4480
rect 2866 4428 2872 4480
rect 2924 4428 2930 4480
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 6288 4468 6316 4508
rect 7285 4505 7297 4508
rect 7331 4505 7343 4539
rect 7285 4499 7343 4505
rect 5307 4440 6316 4468
rect 6733 4471 6791 4477
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 6914 4468 6920 4480
rect 6779 4440 6920 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 6914 4428 6920 4440
rect 6972 4468 6978 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 6972 4440 7205 4468
rect 6972 4428 6978 4440
rect 7193 4437 7205 4440
rect 7239 4468 7251 4471
rect 7834 4468 7840 4480
rect 7239 4440 7840 4468
rect 7239 4437 7251 4440
rect 7193 4431 7251 4437
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 7926 4428 7932 4480
rect 7984 4428 7990 4480
rect 1104 4378 8372 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8372 4378
rect 1104 4304 8372 4326
rect 2038 4224 2044 4276
rect 2096 4264 2102 4276
rect 2096 4236 2774 4264
rect 2096 4224 2102 4236
rect 2130 4156 2136 4208
rect 2188 4196 2194 4208
rect 2654 4199 2712 4205
rect 2654 4196 2666 4199
rect 2188 4168 2666 4196
rect 2188 4156 2194 4168
rect 2654 4165 2666 4168
rect 2700 4165 2712 4199
rect 2746 4196 2774 4236
rect 6086 4224 6092 4276
rect 6144 4224 6150 4276
rect 7742 4224 7748 4276
rect 7800 4224 7806 4276
rect 6914 4196 6920 4208
rect 2746 4168 6920 4196
rect 2654 4159 2712 4165
rect 6914 4156 6920 4168
rect 6972 4156 6978 4208
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 4994 4131 5052 4137
rect 4994 4128 5006 4131
rect 3844 4100 5006 4128
rect 3844 4088 3850 4100
rect 4994 4097 5006 4100
rect 5040 4097 5052 4131
rect 4994 4091 5052 4097
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 6638 4137 6644 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5224 4100 5457 4128
rect 5224 4088 5230 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 6632 4128 6644 4137
rect 6599 4100 6644 4128
rect 5445 4091 5503 4097
rect 6632 4091 6644 4100
rect 6638 4088 6644 4091
rect 6696 4088 6702 4140
rect 1762 4020 1768 4072
rect 1820 4020 1826 4072
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2004 4032 2421 4060
rect 2004 4020 2010 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5316 4032 6377 4060
rect 5316 4020 5322 4032
rect 5460 4004 5488 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 4154 3992 4160 4004
rect 3835 3964 4160 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 5442 3952 5448 4004
rect 5500 3952 5506 4004
rect 2314 3884 2320 3936
rect 2372 3884 2378 3936
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 3510 3924 3516 3936
rect 3200 3896 3516 3924
rect 3200 3884 3206 3896
rect 3510 3884 3516 3896
rect 3568 3924 3574 3936
rect 3881 3927 3939 3933
rect 3881 3924 3893 3927
rect 3568 3896 3893 3924
rect 3568 3884 3574 3896
rect 3881 3893 3893 3896
rect 3927 3893 3939 3927
rect 3881 3887 3939 3893
rect 1104 3834 8372 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 8372 3834
rect 1104 3760 8372 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 3786 3720 3792 3732
rect 1627 3692 3792 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4522 3720 4528 3732
rect 4028 3692 4528 3720
rect 4028 3680 4034 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 4632 3692 5764 3720
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 3418 3652 3424 3664
rect 3375 3624 3424 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 3418 3612 3424 3624
rect 3476 3652 3482 3664
rect 3476 3624 3832 3652
rect 3476 3612 3482 3624
rect 3804 3596 3832 3624
rect 3878 3612 3884 3664
rect 3936 3612 3942 3664
rect 1670 3544 1676 3596
rect 1728 3544 1734 3596
rect 1946 3544 1952 3596
rect 2004 3544 2010 3596
rect 3602 3544 3608 3596
rect 3660 3544 3666 3596
rect 3786 3544 3792 3596
rect 3844 3544 3850 3596
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4632 3584 4660 3692
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5629 3655 5687 3661
rect 5629 3652 5641 3655
rect 5316 3624 5641 3652
rect 5316 3612 5322 3624
rect 5629 3621 5641 3624
rect 5675 3621 5687 3655
rect 5629 3615 5687 3621
rect 4028 3556 4660 3584
rect 4028 3544 4034 3556
rect 1578 3476 1584 3528
rect 1636 3476 1642 3528
rect 1688 3516 1716 3544
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1688 3488 1869 3516
rect 1857 3485 1869 3488
rect 1903 3516 1915 3519
rect 3620 3516 3648 3544
rect 4246 3516 4252 3528
rect 1903 3488 3464 3516
rect 3620 3488 4252 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 2194 3451 2252 3457
rect 2194 3448 2206 3451
rect 1728 3420 2206 3448
rect 1728 3408 1734 3420
rect 2194 3417 2206 3420
rect 2240 3417 2252 3451
rect 2194 3411 2252 3417
rect 3436 3392 3464 3488
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 5350 3516 5356 3528
rect 4387 3488 5356 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5644 3516 5672 3615
rect 5736 3584 5764 3692
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 7837 3655 7895 3661
rect 7837 3652 7849 3655
rect 7432 3624 7849 3652
rect 7432 3612 7438 3624
rect 7837 3621 7849 3624
rect 7883 3621 7895 3655
rect 7837 3615 7895 3621
rect 5736 3556 6316 3584
rect 5902 3516 5908 3528
rect 5644 3488 5908 3516
rect 5902 3476 5908 3488
rect 5960 3516 5966 3528
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 5960 3488 6193 3516
rect 5960 3476 5966 3488
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6288 3516 6316 3556
rect 6437 3519 6495 3525
rect 6437 3516 6449 3519
rect 6288 3488 6449 3516
rect 6181 3479 6239 3485
rect 6437 3485 6449 3488
rect 6483 3485 6495 3519
rect 6437 3479 6495 3485
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 3602 3408 3608 3460
rect 3660 3448 3666 3460
rect 4798 3448 4804 3460
rect 3660 3420 4804 3448
rect 3660 3408 3666 3420
rect 4798 3408 4804 3420
rect 4856 3448 4862 3460
rect 6086 3448 6092 3460
rect 4856 3420 6092 3448
rect 4856 3408 4862 3420
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3380 1823 3383
rect 1854 3380 1860 3392
rect 1811 3352 1860 3380
rect 1811 3349 1823 3352
rect 1765 3343 1823 3349
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 3418 3340 3424 3392
rect 3476 3380 3482 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3476 3352 3801 3380
rect 3476 3340 3482 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 3789 3343 3847 3349
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 5350 3380 5356 3392
rect 4488 3352 5356 3380
rect 4488 3340 4494 3352
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 6822 3380 6828 3392
rect 6420 3352 6828 3380
rect 6420 3340 6426 3352
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7156 3352 7573 3380
rect 7156 3340 7162 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 1104 3290 8372 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8372 3290
rect 1104 3216 8372 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 2222 3176 2228 3188
rect 1627 3148 2228 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 3694 3176 3700 3188
rect 3568 3148 3700 3176
rect 3568 3136 3574 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4154 3176 4160 3188
rect 4019 3148 4160 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4706 3176 4712 3188
rect 4571 3148 4712 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 7098 3176 7104 3188
rect 5368 3148 7104 3176
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 5258 3108 5264 3120
rect 2004 3080 5264 3108
rect 2004 3068 2010 3080
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 2976 3049 3004 3080
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 2694 3043 2752 3049
rect 2694 3040 2706 3043
rect 2372 3012 2706 3040
rect 2372 3000 2378 3012
rect 2694 3009 2706 3012
rect 2740 3009 2752 3043
rect 2694 3003 2752 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3418 3040 3424 3052
rect 3283 3012 3424 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 3694 3000 3700 3052
rect 3752 3000 3758 3052
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3936 3012 4169 3040
rect 3936 3000 3942 3012
rect 4157 3009 4169 3012
rect 4203 3040 4215 3043
rect 5368 3040 5396 3148
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 5442 3068 5448 3120
rect 5500 3068 5506 3120
rect 5920 3080 6408 3108
rect 4203 3012 5396 3040
rect 5460 3040 5488 3068
rect 5920 3052 5948 3080
rect 5638 3043 5696 3049
rect 5638 3040 5650 3043
rect 5460 3012 5650 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 5638 3009 5650 3012
rect 5684 3009 5696 3043
rect 5638 3003 5696 3009
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 6086 3000 6092 3052
rect 6144 3000 6150 3052
rect 6178 3000 6184 3052
rect 6236 3000 6242 3052
rect 6380 3049 6408 3080
rect 6822 3068 6828 3120
rect 6880 3108 6886 3120
rect 7760 3108 7788 3139
rect 6880 3080 7788 3108
rect 6880 3068 6886 3080
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6512 3012 6633 3040
rect 6512 3000 6518 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 6621 3003 6679 3009
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3200 2944 4077 2972
rect 3200 2932 3206 2944
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 4522 2972 4528 2984
rect 4479 2944 4528 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3160 2836 3188 2932
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 3375 2876 5028 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 2832 2808 3188 2836
rect 3237 2839 3295 2845
rect 2832 2796 2838 2808
rect 3237 2805 3249 2839
rect 3283 2836 3295 2839
rect 3970 2836 3976 2848
rect 3283 2808 3976 2836
rect 3283 2805 3295 2808
rect 3237 2799 3295 2805
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 5000 2836 5028 2876
rect 6012 2876 6408 2904
rect 6012 2836 6040 2876
rect 5000 2808 6040 2836
rect 6380 2836 6408 2876
rect 7558 2836 7564 2848
rect 6380 2808 7564 2836
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 1104 2746 8372 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 8372 2746
rect 1104 2672 8372 2694
rect 1670 2592 1676 2644
rect 1728 2592 1734 2644
rect 1762 2592 1768 2644
rect 1820 2632 1826 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 1820 2604 2421 2632
rect 1820 2592 1826 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6454 2632 6460 2644
rect 6227 2604 6460 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6546 2592 6552 2644
rect 6604 2592 6610 2644
rect 7558 2592 7564 2644
rect 7616 2592 7622 2644
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 2332 2536 3801 2564
rect 2332 2505 2360 2536
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 4614 2564 4620 2576
rect 3789 2527 3847 2533
rect 4264 2536 4620 2564
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 2866 2456 2872 2508
rect 2924 2456 2930 2508
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 4264 2505 4292 2536
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 5644 2536 6745 2564
rect 5644 2505 5672 2536
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 7653 2567 7711 2573
rect 7653 2564 7665 2567
rect 6733 2527 6791 2533
rect 6886 2536 7665 2564
rect 4249 2499 4307 2505
rect 3108 2468 4108 2496
rect 3108 2456 3114 2468
rect 2774 2388 2780 2440
rect 2832 2388 2838 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3786 2428 3792 2440
rect 3651 2400 3792 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4080 2360 4108 2468
rect 4249 2465 4261 2499
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 6886 2496 6914 2536
rect 7653 2533 7665 2536
rect 7699 2533 7711 2567
rect 7653 2527 7711 2533
rect 5629 2459 5687 2465
rect 5736 2468 6914 2496
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4448 2360 4476 2459
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5350 2428 5356 2440
rect 4939 2400 5356 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5350 2388 5356 2400
rect 5408 2428 5414 2440
rect 5736 2428 5764 2468
rect 7190 2456 7196 2508
rect 7248 2456 7254 2508
rect 7374 2456 7380 2508
rect 7432 2456 7438 2508
rect 5408 2400 5764 2428
rect 5408 2388 5414 2400
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7156 2400 8033 2428
rect 7156 2388 7162 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 7374 2360 7380 2372
rect 4080 2332 7380 2360
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3421 2295 3479 2301
rect 3421 2292 3433 2295
rect 3292 2264 3433 2292
rect 3292 2252 3298 2264
rect 3421 2261 3433 2264
rect 3467 2261 3479 2295
rect 3421 2255 3479 2261
rect 1104 2202 8372 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8372 2202
rect 1104 2128 8372 2150
<< via1 >>
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 7748 8916 7800 8968
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 2136 8440 2188 8492
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 6184 8508 6236 8560
rect 4712 8440 4764 8492
rect 6092 8483 6144 8492
rect 6092 8449 6101 8483
rect 6101 8449 6135 8483
rect 6135 8449 6144 8483
rect 6092 8440 6144 8449
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 3332 8236 3384 8288
rect 5356 8372 5408 8424
rect 6920 8372 6972 8424
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 4620 8304 4672 8356
rect 5264 8304 5316 8356
rect 6736 8304 6788 8356
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3148 8032 3200 8084
rect 4804 8032 4856 8084
rect 3332 7896 3384 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 2228 7828 2280 7880
rect 4712 7896 4764 7948
rect 5632 7896 5684 7948
rect 7012 8032 7064 8084
rect 6092 7896 6144 7948
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 5908 7828 5960 7880
rect 6644 7871 6696 7880
rect 6644 7837 6678 7871
rect 6678 7837 6696 7871
rect 6644 7828 6696 7837
rect 3240 7692 3292 7744
rect 5448 7692 5500 7744
rect 7104 7692 7156 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1676 7488 1728 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 2596 7463 2648 7472
rect 2596 7429 2614 7463
rect 2614 7429 2648 7463
rect 2596 7420 2648 7429
rect 2872 7420 2924 7472
rect 6092 7463 6144 7472
rect 6092 7429 6101 7463
rect 6101 7429 6135 7463
rect 6135 7429 6144 7463
rect 6092 7420 6144 7429
rect 6736 7420 6788 7472
rect 5356 7352 5408 7404
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 4528 7148 4580 7200
rect 4712 7148 4764 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 5908 6944 5960 6996
rect 3332 6876 3384 6928
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 3240 6740 3292 6792
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 6828 6876 6880 6928
rect 7012 6808 7064 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 6000 6740 6052 6792
rect 7656 6740 7708 6792
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 3056 6672 3108 6724
rect 4712 6672 4764 6724
rect 2136 6604 2188 6656
rect 2596 6604 2648 6656
rect 3608 6604 3660 6656
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 5264 6672 5316 6724
rect 5632 6672 5684 6724
rect 6276 6604 6328 6656
rect 6368 6647 6420 6656
rect 6368 6613 6377 6647
rect 6377 6613 6411 6647
rect 6411 6613 6420 6647
rect 6368 6604 6420 6613
rect 6920 6604 6972 6656
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 4252 6400 4304 6452
rect 5080 6400 5132 6452
rect 5172 6400 5224 6452
rect 5448 6400 5500 6452
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 6092 6400 6144 6452
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 6276 6400 6328 6452
rect 2412 6332 2464 6384
rect 4620 6332 4672 6384
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 2964 6264 3016 6316
rect 3148 6307 3200 6316
rect 3148 6273 3182 6307
rect 3182 6273 3200 6307
rect 3148 6264 3200 6273
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4712 6264 4764 6316
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5448 6264 5500 6316
rect 6460 6332 6512 6384
rect 5632 6264 5684 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 7380 6400 7432 6452
rect 7932 6400 7984 6452
rect 7840 6332 7892 6384
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 4896 6196 4948 6248
rect 6184 6239 6236 6248
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 7104 6196 7156 6248
rect 3240 6060 3292 6112
rect 3976 6060 4028 6112
rect 5264 6060 5316 6112
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 5908 6060 5960 6112
rect 6644 6060 6696 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2596 5856 2648 5908
rect 2964 5899 3016 5908
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 2780 5788 2832 5840
rect 3148 5856 3200 5908
rect 3884 5899 3936 5908
rect 3884 5865 3893 5899
rect 3893 5865 3927 5899
rect 3927 5865 3936 5899
rect 3884 5856 3936 5865
rect 4896 5856 4948 5908
rect 3516 5788 3568 5840
rect 2320 5720 2372 5772
rect 3608 5763 3660 5772
rect 3608 5729 3617 5763
rect 3617 5729 3651 5763
rect 3651 5729 3660 5763
rect 3608 5720 3660 5729
rect 3976 5788 4028 5840
rect 7104 5856 7156 5908
rect 5080 5788 5132 5840
rect 5908 5788 5960 5840
rect 7840 5856 7892 5908
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2412 5627 2464 5636
rect 2412 5593 2421 5627
rect 2421 5593 2455 5627
rect 2455 5593 2464 5627
rect 2412 5584 2464 5593
rect 2504 5627 2556 5636
rect 2504 5593 2513 5627
rect 2513 5593 2547 5627
rect 2547 5593 2556 5627
rect 2504 5584 2556 5593
rect 2872 5584 2924 5636
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6000 5652 6052 5704
rect 6460 5652 6512 5704
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 5172 5584 5224 5636
rect 5724 5584 5776 5636
rect 6368 5584 6420 5636
rect 7656 5584 7708 5636
rect 3884 5516 3936 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4804 5312 4856 5364
rect 6184 5312 6236 5364
rect 2044 5244 2096 5296
rect 2872 5244 2924 5296
rect 3516 5244 3568 5296
rect 2228 5176 2280 5228
rect 2780 5219 2832 5228
rect 2780 5185 2789 5219
rect 2789 5185 2823 5219
rect 2823 5185 2832 5219
rect 2780 5176 2832 5185
rect 1676 5108 1728 5160
rect 3976 5176 4028 5228
rect 3240 5151 3292 5160
rect 3240 5117 3249 5151
rect 3249 5117 3283 5151
rect 3283 5117 3292 5151
rect 3240 5108 3292 5117
rect 2688 5040 2740 5092
rect 3424 5108 3476 5160
rect 4620 5108 4672 5160
rect 3608 5040 3660 5092
rect 4528 5040 4580 5092
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 3700 4972 3752 5024
rect 4712 4972 4764 5024
rect 5908 5244 5960 5296
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 6368 5108 6420 5160
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 7196 5040 7248 5092
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 6644 4972 6696 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2596 4768 2648 4820
rect 2780 4768 2832 4820
rect 7656 4768 7708 4820
rect 1584 4700 1636 4752
rect 2504 4700 2556 4752
rect 3056 4700 3108 4752
rect 3332 4700 3384 4752
rect 6828 4632 6880 4684
rect 7656 4632 7708 4684
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 4160 4564 4212 4616
rect 3700 4496 3752 4548
rect 5448 4564 5500 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 6092 4496 6144 4548
rect 1860 4428 1912 4480
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 2872 4471 2924 4480
rect 2872 4437 2881 4471
rect 2881 4437 2915 4471
rect 2915 4437 2924 4471
rect 2872 4428 2924 4437
rect 6920 4428 6972 4480
rect 7840 4428 7892 4480
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2044 4224 2096 4276
rect 2136 4156 2188 4208
rect 6092 4267 6144 4276
rect 6092 4233 6101 4267
rect 6101 4233 6135 4267
rect 6135 4233 6144 4267
rect 6092 4224 6144 4233
rect 7748 4267 7800 4276
rect 7748 4233 7757 4267
rect 7757 4233 7791 4267
rect 7791 4233 7800 4267
rect 7748 4224 7800 4233
rect 6920 4156 6972 4208
rect 3792 4088 3844 4140
rect 5172 4088 5224 4140
rect 6644 4131 6696 4140
rect 6644 4097 6678 4131
rect 6678 4097 6696 4131
rect 6644 4088 6696 4097
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 1952 4020 2004 4072
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 4160 3952 4212 4004
rect 5448 3952 5500 4004
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 3148 3884 3200 3936
rect 3516 3884 3568 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3792 3680 3844 3732
rect 3976 3680 4028 3732
rect 4528 3680 4580 3732
rect 3424 3612 3476 3664
rect 3884 3655 3936 3664
rect 3884 3621 3893 3655
rect 3893 3621 3927 3655
rect 3927 3621 3936 3655
rect 3884 3612 3936 3621
rect 1676 3544 1728 3596
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 3608 3544 3660 3596
rect 3792 3544 3844 3596
rect 3976 3544 4028 3596
rect 5264 3612 5316 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 4252 3519 4304 3528
rect 1676 3408 1728 3460
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 5356 3476 5408 3528
rect 7380 3612 7432 3664
rect 5908 3476 5960 3528
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 3608 3408 3660 3460
rect 4804 3408 4856 3460
rect 6092 3408 6144 3460
rect 1860 3340 1912 3392
rect 3424 3340 3476 3392
rect 4436 3340 4488 3392
rect 5356 3340 5408 3392
rect 6368 3340 6420 3392
rect 6828 3340 6880 3392
rect 7104 3340 7156 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 2228 3136 2280 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 3700 3136 3752 3188
rect 4160 3136 4212 3188
rect 4712 3136 4764 3188
rect 1952 3068 2004 3120
rect 2320 3000 2372 3052
rect 5264 3068 5316 3120
rect 3424 3000 3476 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 3884 3000 3936 3052
rect 7104 3136 7156 3188
rect 5448 3068 5500 3120
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 6828 3068 6880 3120
rect 6460 3000 6512 3052
rect 3148 2932 3200 2984
rect 4528 2932 4580 2984
rect 2780 2796 2832 2848
rect 3976 2796 4028 2848
rect 7564 2796 7616 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 1768 2592 1820 2644
rect 6460 2592 6512 2644
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 3056 2499 3108 2508
rect 3056 2465 3065 2499
rect 3065 2465 3099 2499
rect 3099 2465 3108 2499
rect 4620 2524 4672 2576
rect 3056 2456 3108 2465
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 3792 2388 3844 2440
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4528 2388 4580 2440
rect 5356 2388 5408 2440
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 7380 2499 7432 2508
rect 7380 2465 7389 2499
rect 7389 2465 7423 2499
rect 7423 2465 7432 2499
rect 7380 2456 7432 2465
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7380 2320 7432 2372
rect 3240 2252 3292 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 7585 1532 8298
rect 1688 7886 1716 8434
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1490 7576 1546 7585
rect 1688 7546 1716 7822
rect 1490 7511 1546 7520
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1872 6905 1900 8298
rect 1858 6896 1914 6905
rect 1858 6831 1914 6840
rect 2148 6662 2176 8434
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6322 2176 6598
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2240 5710 2268 7822
rect 2608 7478 2636 8230
rect 3160 8090 3188 8366
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3344 7954 3372 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 1596 3534 1624 4694
rect 1688 4554 1716 5102
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1688 3602 1716 4490
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 2650 1716 3402
rect 1780 2650 1808 4014
rect 1872 3398 1900 4422
rect 2056 4282 2084 5238
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2240 4622 2268 5170
rect 2332 5030 2360 5714
rect 2424 5642 2452 6326
rect 2608 5914 2636 6598
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2780 5840 2832 5846
rect 2884 5794 2912 7414
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2976 6866 3004 7278
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 6322 3004 6802
rect 3252 6798 3280 7686
rect 3344 6934 3372 7890
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7206 4568 7822
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2964 5908 3016 5914
rect 3068 5896 3096 6666
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3160 5914 3188 6258
rect 3252 6118 3280 6734
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3016 5868 3096 5896
rect 3148 5908 3200 5914
rect 2964 5850 3016 5856
rect 3148 5850 3200 5856
rect 2832 5788 2912 5794
rect 2780 5782 2912 5788
rect 2792 5766 2912 5782
rect 3238 5808 3294 5817
rect 3238 5743 3294 5752
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2516 4758 2544 5578
rect 2884 5302 2912 5578
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4826 2636 4966
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2148 4214 2176 4422
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1964 3602 1992 4014
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1964 3126 1992 3538
rect 2240 3194 2268 4558
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 2332 3058 2360 3878
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2700 2530 2728 5034
rect 2792 4826 2820 5170
rect 3252 5166 3280 5743
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3344 4758 3372 6870
rect 3608 6792 3660 6798
rect 3528 6752 3608 6780
rect 3528 6361 3556 6752
rect 3608 6734 3660 6740
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 3514 6352 3570 6361
rect 3514 6287 3570 6296
rect 3528 5846 3556 6287
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3620 5778 3648 6598
rect 4264 6458 4292 6598
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4632 6390 4660 8298
rect 4724 7954 4752 8434
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 8090 4844 8230
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6730 4752 7142
rect 5276 6730 5304 8298
rect 5368 7886 5396 8366
rect 6104 7954 6132 8434
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 5356 7880 5408 7886
rect 5408 7840 5580 7868
rect 5356 7822 5408 7828
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4066 6216 4122 6225
rect 4540 6202 4568 6258
rect 4540 6174 4660 6202
rect 4066 6151 4122 6160
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3896 5574 3924 5850
rect 3988 5846 4016 6054
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4080 5710 4108 6151
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2608 2502 2728 2530
rect 2608 800 2636 2502
rect 2792 2446 2820 2790
rect 2884 2514 2912 4422
rect 3068 2514 3096 4694
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 2990 3188 3878
rect 3436 3670 3464 5102
rect 3528 4622 3556 5238
rect 3988 5234 4016 5646
rect 4632 5250 4660 6174
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4540 5222 4660 5250
rect 4724 5250 4752 6258
rect 4804 6248 4856 6254
rect 4802 6216 4804 6225
rect 4896 6248 4948 6254
rect 4856 6216 4858 6225
rect 4896 6190 4948 6196
rect 4802 6151 4858 6160
rect 4816 5370 4844 6151
rect 4908 5914 4936 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5817 5028 6258
rect 5092 5846 5120 6394
rect 5080 5840 5132 5846
rect 4986 5808 5042 5817
rect 5080 5782 5132 5788
rect 4986 5743 5042 5752
rect 5184 5642 5212 6394
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4724 5222 4844 5250
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3528 3942 3556 4558
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3424 3664 3476 3670
rect 3620 3618 3648 5034
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3712 4554 3740 4966
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3804 3738 3832 4082
rect 3988 3738 4016 5170
rect 4540 5098 4568 5222
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4172 4026 4200 4558
rect 4080 4010 4200 4026
rect 4080 4004 4212 4010
rect 4080 3998 4160 4004
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3424 3606 3476 3612
rect 3528 3602 3648 3618
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 4080 3618 4108 3998
rect 4160 3946 4212 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 3528 3596 3660 3602
rect 3528 3590 3608 3596
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 3058 3464 3334
rect 3528 3194 3556 3590
rect 3608 3538 3660 3544
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3620 3058 3648 3402
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3712 3058 3740 3130
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3804 2446 3832 3538
rect 3896 3058 3924 3606
rect 3976 3596 4028 3602
rect 4080 3590 4200 3618
rect 3976 3538 4028 3544
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3988 2854 4016 3538
rect 4172 3194 4200 3590
rect 4252 3528 4304 3534
rect 4304 3476 4476 3482
rect 4252 3470 4476 3476
rect 4264 3454 4476 3470
rect 4448 3398 4476 3454
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4172 2938 4200 3130
rect 4540 2990 4568 3674
rect 4080 2910 4200 2938
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 4080 2530 4108 2910
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2582 4660 5102
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 3194 4752 4966
rect 4816 3466 4844 5222
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5276 4162 5304 6054
rect 5368 5574 5396 7346
rect 5460 6458 5488 7686
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5552 6361 5580 7840
rect 5644 6730 5672 7890
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7002 5948 7822
rect 6104 7478 6132 7890
rect 6092 7472 6144 7478
rect 6012 7432 6092 7460
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6012 6798 6040 7432
rect 6092 7414 6144 7420
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5538 6352 5594 6361
rect 5448 6316 5500 6322
rect 5644 6322 5672 6666
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5538 6287 5594 6296
rect 5632 6316 5684 6322
rect 5448 6258 5500 6264
rect 5632 6258 5684 6264
rect 5460 6225 5488 6258
rect 5446 6216 5502 6225
rect 5446 6151 5502 6160
rect 5920 6118 5948 6394
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5736 5642 5764 6054
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5184 4146 5304 4162
rect 5172 4140 5304 4146
rect 5224 4134 5304 4140
rect 5172 4082 5224 4088
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3670 5304 4014
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5276 3126 5304 3606
rect 5368 3534 5396 5510
rect 5920 5302 5948 5782
rect 6012 5710 6040 6734
rect 6196 6458 6224 8502
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7886 6684 8230
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6748 7478 6776 8298
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6828 6928 6880 6934
rect 6366 6896 6422 6905
rect 6828 6870 6880 6876
rect 6366 6831 6422 6840
rect 6380 6662 6408 6831
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6288 6458 6316 6598
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6104 6361 6132 6394
rect 6460 6384 6512 6390
rect 6090 6352 6146 6361
rect 6460 6326 6512 6332
rect 6550 6352 6606 6361
rect 6090 6287 6146 6296
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6196 5370 6224 6190
rect 6380 5642 6408 6258
rect 6472 5710 6500 6326
rect 6550 6287 6552 6296
rect 6604 6287 6606 6296
rect 6644 6316 6696 6322
rect 6552 6258 6604 6264
rect 6644 6258 6696 6264
rect 6656 6118 6684 6258
rect 6840 6254 6868 6870
rect 6932 6662 6960 8366
rect 7024 8090 7052 8910
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 6866 7144 7686
rect 7208 7585 7236 8774
rect 7194 7576 7250 7585
rect 7194 7511 7250 7520
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7024 6662 7052 6802
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6840 5817 6868 6190
rect 6826 5808 6882 5817
rect 6826 5743 6882 5752
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4010 5488 4558
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6104 4282 6132 4490
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5368 3074 5396 3334
rect 5448 3120 5500 3126
rect 5368 3068 5448 3074
rect 5368 3062 5500 3068
rect 5368 3046 5488 3062
rect 5920 3058 5948 3470
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6104 3058 6132 3402
rect 6196 3058 6224 4966
rect 6380 3398 6408 5102
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4146 6684 4966
rect 6840 4690 6868 5743
rect 7024 5234 7052 6598
rect 7392 6458 7420 8774
rect 7760 7546 7788 8910
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7760 6882 7788 7482
rect 7668 6854 7788 6882
rect 7668 6798 7696 6854
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7760 6644 7788 6734
rect 7668 6616 7788 6644
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 5914 7144 6190
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7668 5642 7696 6616
rect 7852 6390 7880 6734
rect 7944 6458 7972 8366
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7852 5914 7880 6326
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7668 5250 7696 5578
rect 7668 5234 7880 5250
rect 8036 5234 8064 5646
rect 7012 5228 7064 5234
rect 7668 5228 7892 5234
rect 7668 5222 7840 5228
rect 7012 5170 7064 5176
rect 7840 5170 7892 5176
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4214 6960 4422
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6550 3496 6606 3505
rect 6550 3431 6606 3440
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 5908 3052 5960 3058
rect 4620 2576 4672 2582
rect 4080 2502 4200 2530
rect 4620 2518 4672 2524
rect 4172 2446 4200 2502
rect 5368 2446 5396 3046
rect 5908 2994 5960 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6380 2446 6408 3334
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6472 2650 6500 2994
rect 6564 2650 6592 3431
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6840 3126 6868 3334
rect 7116 3194 7144 3334
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 7116 2446 7144 3130
rect 7208 2514 7236 5034
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7392 2514 7420 3606
rect 7668 3534 7696 4626
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7760 4282 7788 4558
rect 7852 4486 7880 5170
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7944 4185 7972 4422
rect 7930 4176 7986 4185
rect 7930 4111 7986 4120
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7576 2650 7604 2790
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 800 3280 2246
rect 4540 800 4568 2382
rect 7392 2378 7420 2450
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
<< via2 >>
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 1490 7520 1546 7576
rect 1858 6840 1914 6896
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3238 5752 3294 5808
rect 3514 6296 3570 6352
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4066 6160 4122 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4802 6196 4804 6216
rect 4804 6196 4856 6216
rect 4856 6196 4858 6216
rect 4802 6160 4858 6196
rect 4986 5752 5042 5808
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 5538 6296 5594 6352
rect 5446 6160 5502 6216
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 6366 6840 6422 6896
rect 6090 6296 6146 6352
rect 6550 6316 6606 6352
rect 6550 6296 6552 6316
rect 6552 6296 6604 6316
rect 6604 6296 6606 6316
rect 7194 7520 7250 7576
rect 6826 5752 6882 5808
rect 6550 3440 6606 3496
rect 7930 4120 7986 4176
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 7189 7578 7255 7581
rect 8746 7578 9546 7608
rect 7189 7576 9546 7578
rect 7189 7520 7194 7576
rect 7250 7520 9546 7576
rect 7189 7518 9546 7520
rect 7189 7515 7255 7518
rect 8746 7488 9546 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 1853 6898 1919 6901
rect 0 6896 1919 6898
rect 0 6840 1858 6896
rect 1914 6840 1919 6896
rect 0 6838 1919 6840
rect 0 6808 800 6838
rect 1853 6835 1919 6838
rect 6361 6898 6427 6901
rect 8746 6898 9546 6928
rect 6361 6896 9546 6898
rect 6361 6840 6366 6896
rect 6422 6840 9546 6896
rect 6361 6838 9546 6840
rect 6361 6835 6427 6838
rect 8746 6808 9546 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 3509 6354 3575 6357
rect 5533 6354 5599 6357
rect 6085 6354 6151 6357
rect 6545 6354 6611 6357
rect 3509 6352 6611 6354
rect 3509 6296 3514 6352
rect 3570 6296 5538 6352
rect 5594 6296 6090 6352
rect 6146 6296 6550 6352
rect 6606 6296 6611 6352
rect 3509 6294 6611 6296
rect 3509 6291 3575 6294
rect 5533 6291 5599 6294
rect 6085 6291 6151 6294
rect 6545 6291 6611 6294
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 4797 6218 4863 6221
rect 5441 6218 5507 6221
rect 4797 6216 5507 6218
rect 4797 6160 4802 6216
rect 4858 6160 5446 6216
rect 5502 6160 5507 6216
rect 4797 6158 5507 6160
rect 4797 6155 4863 6158
rect 5441 6155 5507 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 3233 5810 3299 5813
rect 4981 5810 5047 5813
rect 6821 5810 6887 5813
rect 3233 5808 6887 5810
rect 3233 5752 3238 5808
rect 3294 5752 4986 5808
rect 5042 5752 6826 5808
rect 6882 5752 6887 5808
rect 3233 5750 6887 5752
rect 3233 5747 3299 5750
rect 4981 5747 5047 5750
rect 6821 5747 6887 5750
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 7925 4178 7991 4181
rect 8746 4178 9546 4208
rect 7925 4176 9546 4178
rect 7925 4120 7930 4176
rect 7986 4120 9546 4176
rect 7925 4118 9546 4120
rect 7925 4115 7991 4118
rect 8746 4088 9546 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 6545 3498 6611 3501
rect 8746 3498 9546 3528
rect 6545 3496 9546 3498
rect 6545 3440 6550 3496
rect 6606 3440 9546 3496
rect 6545 3438 9546 3440
rect 6545 3435 6611 3438
rect 8746 3408 9546 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9296
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9296
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _34_
timestamp -3599
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _35_
timestamp -3599
transform -1 0 3772 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _36_
timestamp -3599
transform 1 0 6716 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _37_
timestamp -3599
transform 1 0 2392 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _38_
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _39_
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _40_
timestamp -3599
transform 1 0 2392 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _41_
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _42_
timestamp -3599
transform -1 0 7544 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _43_
timestamp -3599
transform 1 0 6624 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _44_
timestamp -3599
transform -1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _45_
timestamp -3599
transform -1 0 4324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _46_
timestamp -3599
transform -1 0 3680 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _47_
timestamp -3599
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _48_
timestamp -3599
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _49_
timestamp -3599
transform 1 0 2576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _50_
timestamp -3599
transform 1 0 3680 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _51_
timestamp -3599
transform -1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _52_
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _53_
timestamp -3599
transform -1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _54_
timestamp -3599
transform -1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _55_
timestamp -3599
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _56_
timestamp -3599
transform -1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _57_
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _58_
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _59_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _60_
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _61_
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _62_
timestamp -3599
transform -1 0 8004 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _63_
timestamp -3599
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _64_
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _65_
timestamp -3599
transform 1 0 4968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _66_
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _67_
timestamp -3599
transform 1 0 4600 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _68_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _69_
timestamp -3599
transform -1 0 3036 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _70_
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _71_
timestamp -3599
transform -1 0 3036 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _72_
timestamp -3599
transform -1 0 2944 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _73_
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _74_
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _75_
timestamp -3599
transform 1 0 6348 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _76_
timestamp -3599
transform 1 0 6164 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _77_
timestamp -3599
transform -1 0 5336 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _78_
timestamp -3599
transform 1 0 2392 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _79_
timestamp -3599
transform 1 0 2944 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _80_
timestamp -3599
transform 1 0 2852 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _81_
timestamp -3599
transform 1 0 5336 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _82_
timestamp -3599
transform 1 0 5888 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _83_
timestamp -3599
transform 1 0 4784 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _84_
timestamp -3599
transform -1 0 5980 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_21
timestamp -3599
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_73
timestamp -3599
transform 1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp -3599
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp -3599
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_46
timestamp -3599
transform 1 0 5336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_73
timestamp -3599
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp -3599
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp -3599
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp -3599
transform 1 0 7452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp -3599
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_73
timestamp -3599
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp -3599
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_39
timestamp -3599
transform 1 0 4692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_73
timestamp -3599
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp -3599
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_24
timestamp -3599
transform 1 0 3312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_32
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_43
timestamp -3599
transform 1 0 5060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp -3599
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636964856
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636964856
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -3599
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636964856
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636964856
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_53
timestamp -3599
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_57
timestamp -3599
transform 1 0 6348 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_63
timestamp -3599
transform 1 0 6900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -3599
transform -1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -3599
transform 1 0 4784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -3599
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -3599
transform -1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -3599
transform 1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -3599
transform -1 0 2392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -3599
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -3599
transform -1 0 3680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp -3599
transform -1 0 4692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp -3599
transform -1 0 3680 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp -3599
transform 1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp -3599
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp -3599
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform -1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform -1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_30
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_31
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_32
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_34
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_35
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_36
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_37
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_38
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_39
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_40
timestamp -3599
transform 1 0 6256 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 analog_out
port 2 nsew signal input
flabel metal3 s 8746 3408 9546 3528 0 FreeSans 480 0 0 0 b[0]
port 3 nsew signal output
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 b[1]
port 4 nsew signal output
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 b[2]
port 5 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 b[3]
port 6 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 b[4]
port 7 nsew signal output
flabel metal3 s 8746 4088 9546 4208 0 FreeSans 480 0 0 0 b[5]
port 8 nsew signal output
flabel metal3 s 8746 6808 9546 6928 0 FreeSans 480 0 0 0 b[6]
port 9 nsew signal output
flabel metal3 s 8746 7488 9546 7608 0 FreeSans 480 0 0 0 b[7]
port 10 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 clk
port 11 nsew signal input
rlabel metal1 4738 8704 4738 8704 0 VGND
rlabel metal1 4738 9248 4738 9248 0 VPWR
rlabel metal1 5658 2516 5658 2516 0 _00_
rlabel metal1 2116 2618 2116 2618 0 _01_
rlabel metal1 2346 2516 2346 2516 0 _02_
rlabel metal2 3634 6188 3634 6188 0 _03_
rlabel metal2 3174 8228 3174 8228 0 _04_
rlabel metal1 7268 4794 7268 4794 0 _05_
rlabel metal1 7728 6426 7728 6426 0 _06_
rlabel metal1 6808 6630 6808 6630 0 _07_
rlabel metal1 3634 2822 3634 2822 0 _08_
rlabel metal2 3818 3910 3818 3910 0 _09_
rlabel metal1 2422 4182 2422 4182 0 _10_
rlabel via1 2806 5797 2806 5797 0 _11_
rlabel metal1 2990 5814 2990 5814 0 _12_
rlabel metal1 5336 4114 5336 4114 0 _13_
rlabel metal1 5964 5610 5964 5610 0 _14_
rlabel metal1 5193 6698 5193 6698 0 _15_
rlabel metal2 3634 3230 3634 3230 0 _16_
rlabel metal2 5014 6035 5014 6035 0 _17_
rlabel metal1 6992 2822 6992 2822 0 _18_
rlabel metal1 1794 3502 1794 3502 0 _19_
rlabel metal2 1610 4114 1610 4114 0 _20_
rlabel metal1 2300 4794 2300 4794 0 _21_
rlabel metal1 4370 5202 4370 5202 0 _22_
rlabel metal2 3726 4760 3726 4760 0 _23_
rlabel metal2 2438 5984 2438 5984 0 _24_
rlabel metal1 2668 5882 2668 5882 0 _25_
rlabel metal1 3818 5644 3818 5644 0 _26_
rlabel metal1 4416 5882 4416 5882 0 _27_
rlabel metal1 5566 6154 5566 6154 0 _28_
rlabel metal2 4830 5780 4830 5780 0 _29_
rlabel metal1 5750 6290 5750 6290 0 _30_
rlabel metal1 6946 5270 6946 5270 0 _31_
rlabel metal1 4922 8058 4922 8058 0 _32_
rlabel metal1 5536 8534 5536 8534 0 _33_
rlabel metal2 4554 1588 4554 1588 0 analog_out
rlabel metal3 7736 3468 7736 3468 0 b[0]
rlabel metal2 2622 1639 2622 1639 0 b[1]
rlabel metal2 3266 1520 3266 1520 0 b[2]
rlabel metal3 1280 6868 1280 6868 0 b[3]
rlabel metal3 1096 7548 1096 7548 0 b[4]
rlabel metal2 7958 4301 7958 4301 0 b[5]
rlabel metal2 6394 6749 6394 6749 0 b[6]
rlabel metal2 7222 8177 7222 8177 0 b[7]
rlabel metal2 4094 5933 4094 5933 0 clk
rlabel metal2 5382 4522 5382 4522 0 clknet_0_clk
rlabel metal1 2208 4046 2208 4046 0 clknet_1_0__leaf_clk
rlabel metal1 6256 7922 6256 7922 0 clknet_1_1__leaf_clk
rlabel metal1 7590 2414 7590 2414 0 counter\[0\]
rlabel metal1 3634 2958 3634 2958 0 counter\[1\]
rlabel metal2 4186 2465 4186 2465 0 counter\[2\]
rlabel metal1 4554 6698 4554 6698 0 counter\[3\]
rlabel metal1 4140 6086 4140 6086 0 counter\[4\]
rlabel metal1 2116 5270 2116 5270 0 counter\[5\]
rlabel metal1 7498 6358 7498 6358 0 counter\[6\]
rlabel metal1 6072 6970 6072 6970 0 counter\[7\]
rlabel metal1 7291 2550 7291 2550 0 net1
rlabel metal2 7406 2414 7406 2414 0 net10
rlabel metal1 6808 4522 6808 4522 0 net11
rlabel via1 6665 4114 6665 4114 0 net12
rlabel metal1 6348 5066 6348 5066 0 net13
rlabel metal1 6348 2618 6348 2618 0 net14
rlabel metal1 2622 7786 2622 7786 0 net15
rlabel via1 2626 7446 2626 7446 0 net16
rlabel metal2 2898 3468 2898 3468 0 net17
rlabel metal1 2534 3026 2534 3026 0 net18
rlabel metal1 7222 6426 7222 6426 0 net19
rlabel metal1 5658 5134 5658 5134 0 net2
rlabel metal1 6711 7446 6711 7446 0 net20
rlabel metal2 7130 7276 7130 7276 0 net21
rlabel via1 6665 7854 6665 7854 0 net22
rlabel metal1 4278 2516 4278 2516 0 net23
rlabel metal2 1702 3026 1702 3026 0 net24
rlabel metal1 3542 6426 3542 6426 0 net25
rlabel metal2 3036 5882 3036 5882 0 net26
rlabel metal2 6210 4012 6210 4012 0 net27
rlabel metal2 6118 4386 6118 4386 0 net28
rlabel metal1 3128 7854 3128 7854 0 net29
rlabel metal2 2254 3876 2254 3876 0 net3
rlabel metal1 1702 4454 1702 4454 0 net30
rlabel metal1 7268 5678 7268 5678 0 net31
rlabel metal1 6302 5338 6302 5338 0 net32
rlabel metal2 2806 4998 2806 4998 0 net33
rlabel metal1 3726 2414 3726 2414 0 net4
rlabel metal1 1886 6630 1886 6630 0 net5
rlabel metal2 1702 7684 1702 7684 0 net6
rlabel metal1 6670 4590 6670 4590 0 net7
rlabel metal2 7774 8228 7774 8228 0 net8
rlabel metal1 6762 8058 6762 8058 0 net9
rlabel metal1 3772 5202 3772 5202 0 out_d
<< properties >>
string FIXED_BBOX 0 0 9546 11690
<< end >>
