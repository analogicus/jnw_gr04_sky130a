magic
tech sky130A
magscale 1 2
timestamp 1744566163
<< locali >>
rect -5108 7250 -4444 7258
rect -5108 7070 -4974 7250
rect -4794 7070 -4444 7250
rect -5108 7066 -4444 7070
rect -2316 7066 -1808 7258
rect -2048 6868 -1808 7066
rect -2048 6688 -2002 6868
rect -1822 6688 -1808 6868
rect -2048 6168 -1808 6688
rect -2048 6106 -1986 6168
rect -2619 6012 -1986 6106
rect -1830 6106 -1808 6168
rect -1830 6012 -1743 6106
rect -2619 5728 -1743 6012
rect 2518 2573 3434 2717
rect -2702 1690 -2510 1718
rect -2702 1360 -2510 1578
rect -1550 1420 -1256 1745
rect -1550 1360 3987 1420
rect -4678 1304 3987 1360
rect -4678 1249 -1252 1304
rect -4678 236 -1230 1249
rect -274 1152 -200 1155
rect -274 1150 -204 1152
rect -274 1088 -208 1150
rect -274 1083 -199 1088
rect -4678 204 -1165 236
rect -4679 170 -1165 204
rect -4679 139 -1261 170
rect -4679 129 -1165 139
rect -1101 129 -1029 265
rect 3871 129 3987 1304
rect -4679 105 5169 129
rect -4678 40 5169 105
rect -1411 30 5169 40
rect -1371 -265 -1165 30
<< viali >>
rect -4974 7070 -4794 7250
rect -2002 6688 -1822 6868
rect -3190 6348 -3138 6400
rect 358 6544 410 6596
rect -1986 6012 -1830 6168
rect 434 3167 488 3221
rect 994 2371 1038 2427
rect 1492 2377 1536 2421
rect 2377 2371 2437 2443
rect 2778 2377 2838 2437
rect 3660 2371 3720 2443
rect 4062 2377 4122 2437
rect 187 1481 259 1541
rect 4051 1481 4123 1541
rect -199 1083 -139 1155
rect 196 1089 256 1149
rect 1080 1089 1140 1149
rect 1482 1083 1542 1155
rect 2354 1089 2414 1149
rect 2763 1083 2823 1155
rect 3665 1083 3725 1155
rect 4057 1086 4117 1146
<< metal1 >>
rect -2702 7460 -2510 7466
rect -2880 7268 -2702 7460
rect -4980 7250 -4788 7262
rect -4980 7070 -4974 7250
rect -4794 7070 -4788 7250
rect -4980 6874 -4788 7070
rect -3942 6938 -2860 7002
rect -2830 6938 -2766 7268
rect -2702 7262 -2510 7268
rect -4980 6682 -4254 6874
rect -4132 6682 -2576 6874
rect -2508 6868 -1810 6874
rect -2508 6688 -2002 6868
rect -1822 6688 -1810 6868
rect -2508 6682 -1810 6688
rect 346 6538 352 6602
rect 416 6538 422 6602
rect -4878 6296 -4366 6488
rect -3196 6400 -3132 6412
rect -3196 6348 -3190 6400
rect -3138 6348 -3132 6400
rect -3196 6312 -3132 6348
rect -2264 6368 -2200 6374
rect -3202 6248 -3196 6312
rect -3132 6248 -3126 6312
rect -2264 6298 -2200 6304
rect -1998 6168 -1690 6174
rect -1998 6012 -1986 6168
rect -1830 6012 -1690 6168
rect -1998 6006 -1690 6012
rect -1230 6172 -1062 6178
rect -1230 5998 -1062 6004
rect -1680 4360 -1616 4366
rect -682 4362 -490 4368
rect -1680 4290 -1616 4296
rect -1192 4356 -1128 4362
rect -1192 4286 -1128 4292
rect -682 4164 -490 4170
rect -1192 3642 -1128 3682
rect -1192 3538 -1128 3578
rect 422 3221 500 3227
rect 422 3167 434 3221
rect 488 3167 500 3221
rect 422 3161 500 3167
rect 175 1541 271 1547
rect 175 1481 187 1541
rect 259 1481 271 1541
rect 175 1475 271 1481
rect -205 1155 -133 1167
rect 187 1155 259 1475
rect -205 1083 -199 1155
rect -139 1149 268 1155
rect -139 1089 196 1149
rect 256 1089 268 1149
rect -139 1083 268 1089
rect -205 1071 -133 1083
rect -862 958 -798 964
rect -916 952 -862 958
rect 428 949 494 3161
rect 2371 2443 2443 2455
rect 3654 2443 3726 2455
rect 4056 2443 4128 2449
rect 988 2427 1044 2439
rect 1486 2427 1542 2433
rect 988 2371 994 2427
rect 1038 2421 1542 2427
rect 1038 2377 1492 2421
rect 1536 2377 1542 2421
rect 1038 2371 1542 2377
rect 988 2359 1044 2371
rect 1486 2365 1542 2371
rect 2371 2371 2377 2443
rect 2437 2437 2850 2443
rect 2437 2377 2778 2437
rect 2838 2377 2850 2437
rect 2437 2371 2850 2377
rect 3654 2371 3660 2443
rect 3720 2437 4128 2443
rect 3720 2377 4062 2437
rect 4122 2377 4128 2437
rect 3720 2371 4128 2377
rect 2371 2359 2443 2371
rect 3654 2359 3726 2371
rect 4056 2365 4128 2371
rect 907 2122 4293 2188
rect 4039 1541 4135 1547
rect 4039 1481 4051 1541
rect 4123 1481 4135 1541
rect 4039 1475 4135 1481
rect 1476 1155 1548 1167
rect 2757 1155 2829 1167
rect 1068 1149 1482 1155
rect 1068 1089 1080 1149
rect 1140 1089 1482 1149
rect 1068 1083 1482 1089
rect 1542 1083 1548 1155
rect 2342 1149 2763 1155
rect 2342 1089 2354 1149
rect 2414 1089 2763 1149
rect 2342 1083 2763 1089
rect 2823 1083 2829 1155
rect 1476 1071 1548 1083
rect 2757 1071 2829 1083
rect 3659 1155 3731 1167
rect 4051 1155 4123 1475
rect 3659 1083 3665 1155
rect 3725 1146 4124 1155
rect 3725 1086 4057 1146
rect 4117 1086 4124 1146
rect 3725 1083 4124 1086
rect 3659 1071 3731 1083
rect 4051 1074 4123 1083
rect 4292 949 4358 1719
rect -862 888 -798 894
rect -916 882 -798 888
rect 407 883 4358 949
rect -862 842 -798 882
<< via1 >>
rect -2702 7268 -2510 7460
rect 352 6596 416 6602
rect 352 6544 358 6596
rect 358 6544 410 6596
rect 410 6544 416 6596
rect 352 6538 416 6544
rect -3196 6248 -3132 6312
rect -2264 6304 -2200 6368
rect -1230 6004 -1062 6172
rect -1680 4296 -1616 4360
rect -1192 4292 -1128 4356
rect -682 4170 -490 4362
rect -1192 3578 -1128 3642
rect -862 894 -798 958
<< metal2 >>
rect -2507 7460 -2325 7464
rect -2708 7268 -2702 7460
rect -2510 7455 -2320 7460
rect -2510 7273 -2507 7455
rect -2325 7273 -2320 7455
rect -2510 7268 -2320 7273
rect -2507 7264 -2325 7268
rect 352 6602 416 6608
rect -1680 6538 352 6602
rect -1680 6368 -1616 6538
rect 352 6532 416 6538
rect -3196 6312 -3132 6318
rect -2270 6304 -2264 6368
rect -2200 6304 -1616 6368
rect -3196 6168 -3132 6248
rect -3201 6112 -3192 6168
rect -3136 6112 -3127 6168
rect -3196 6108 -3132 6112
rect -1680 4360 -1616 6304
rect -1230 6286 -1062 6295
rect -1236 6004 -1230 6172
rect -1062 6004 -1056 6172
rect -1201 5642 -1192 5706
rect -1136 5642 -1127 5706
rect -1686 4296 -1680 4360
rect -1616 4296 -1610 4360
rect -1192 4356 -1128 5642
rect -682 4480 -490 4489
rect -1198 4292 -1192 4356
rect -1128 4292 -1122 4356
rect -688 4170 -682 4362
rect -490 4170 -484 4362
rect -1198 3578 -1192 3642
rect -1128 3578 -1122 3642
rect -1192 958 -1128 3578
rect -1192 894 -862 958
rect -798 894 -792 958
<< via2 >>
rect -2507 7273 -2325 7455
rect -3192 6112 -3136 6168
rect -1230 6172 -1062 6286
rect -1230 6128 -1062 6172
rect -1192 5642 -1136 5706
rect -682 4362 -490 4480
rect -682 4298 -490 4362
<< metal3 >>
rect -2245 7460 -2055 7465
rect -2512 7459 -2054 7460
rect -2512 7455 -2245 7459
rect -2512 7273 -2507 7455
rect -2325 7273 -2245 7455
rect -2512 7269 -2245 7273
rect -2055 7269 -2054 7459
rect -2512 7268 -2054 7269
rect -2245 7263 -2055 7268
rect -1230 6291 -1062 6800
rect -1235 6286 -1057 6291
rect -3196 6173 -3132 6186
rect -3197 6168 -3131 6173
rect -3197 6112 -3192 6168
rect -3136 6112 -3131 6168
rect -1235 6128 -1230 6286
rect -1062 6128 -1057 6286
rect -1235 6123 -1057 6128
rect -3197 6107 -3131 6112
rect -3196 5706 -3132 6107
rect -1197 5706 -1131 5711
rect -3196 5642 -1192 5706
rect -1136 5642 -1131 5706
rect -1197 5637 -1131 5642
rect -682 4600 -490 4606
rect -687 4298 -682 4485
rect -490 4298 -485 4485
rect -687 4293 -485 4298
<< via3 >>
rect -2245 7269 -2055 7459
rect -682 4480 -490 4600
rect -682 4410 -490 4480
<< metal4 >>
rect -2246 7459 -1826 7460
rect -2246 7269 -2245 7459
rect -2055 7269 -1826 7459
rect -1700 7416 -1572 7476
rect -2246 7268 -1826 7269
rect -2018 6582 -1826 7268
rect -1702 6700 -1580 6760
rect -868 6582 -676 6800
rect -2018 6390 -490 6582
rect -682 4601 -490 6390
rect -683 4600 -489 4601
rect -683 4410 -682 4600
rect -490 4410 -489 4600
rect -683 4409 -489 4410
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1737662937
transform 1 0 3862 0 1 1292
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1737662937
transform 1 0 2574 0 1 1292
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1737662937
transform 1 0 3862 0 1 4
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1737662937
transform 1 0 2574 0 1 4
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1737662937
transform 1 0 -2 0 1 1292
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1737662937
transform 1 0 1286 0 1 1292
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1737662937
transform 1 0 1286 0 1 4
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1737662937
transform 1 0 -2 0 1 4
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  xb1
timestamp 1737662937
transform 1 0 -1290 0 1 4
box 0 0 1340 1340
use JNWTR_CAPX1  xc1 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 -1700 0 1 6700
box 0 0 1080 1080
use JNWATR_PCH_4C5F0  xm4 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 0 1 -3796 -1 0 7162
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xm5
timestamp 1734044400
transform 0 1 -2964 -1 0 7162
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xm6
timestamp 1734044400
transform 0 1 -4596 -1 0 7162
box -184 -128 1336 928
use Opamp_test  xo1
timestamp 1744566163
transform 1 0 -6922 0 1 -246
box 2222 1594 6906 6420
use JNWTR_RPPO16  xr1 ../JNW_TR_SKY130A
timestamp 1744547463
transform 0 -1 3450 -1 0 7061
box 0 0 4472 3440
<< labels >>
flabel metal1 -4878 6296 -4366 6488 0 FreeSans 1600 0 0 0 I_out
port 1 nsew
flabel locali -5108 7066 -4916 7258 0 FreeSans 1600 0 0 0 VDD_1V8
port 2 nsew
flabel locali -1371 -265 -1261 236 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
<< end >>
