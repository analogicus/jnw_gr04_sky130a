magic
tech sky130A
magscale 1 2
timestamp 1744227397
<< locali >>
rect -292 2488 -52 3066
rect -292 2332 -250 2488
rect -94 2332 -52 2488
rect -292 2008 -52 2332
rect 940 2038 1132 3098
rect 1040 1670 1512 1782
rect -1478 768 -1286 1560
rect -290 666 -49 1608
rect 940 762 1132 1588
rect 2596 1518 2860 1778
rect 2620 1278 2860 1518
rect -1478 -340 -1286 218
rect 940 -262 1132 218
rect -1478 -1290 -1286 -838
rect -326 -1242 -20 -790
rect 940 -1186 1132 -838
rect -292 -1272 -20 -1242
rect -260 -1278 -20 -1272
rect -1478 -2108 -1286 -1806
rect -326 -2108 -20 -1758
rect 940 -2108 1132 -1806
rect -1478 -2110 1132 -2108
rect -1478 -2114 562 -2110
rect -1478 -2294 -1088 -2114
rect -908 -2290 562 -2114
rect 742 -2290 1132 -2110
rect -908 -2294 1132 -2290
rect -1478 -2300 1132 -2294
<< viali >>
rect -250 2332 -94 2488
rect 1754 1306 1806 1358
rect -1088 -2294 -908 -2114
rect 562 -2290 742 -2110
<< metal1 >>
rect -242 2494 356 2498
rect -698 2488 356 2494
rect -698 2332 -250 2488
rect -94 2332 356 2488
rect -698 2330 356 2332
rect -698 2326 -82 2330
rect -698 2000 -530 2326
rect 188 2000 356 2330
rect -1094 1102 -902 1640
rect 44 1572 108 1578
rect -460 1508 -454 1572
rect -390 1508 -384 1572
rect 44 1364 108 1508
rect 556 1364 748 1776
rect 44 1358 1818 1364
rect 44 1306 1754 1358
rect 1806 1306 1818 1358
rect 44 1300 1818 1306
rect 400 1236 464 1242
rect -826 1228 -762 1234
rect -762 1164 -390 1228
rect -826 1158 -762 1164
rect -1094 1100 -522 1102
rect -1094 932 -700 1100
rect -532 932 -518 1100
rect -1094 928 -518 932
rect -1094 910 -522 928
rect -698 658 -530 910
rect -454 762 -390 1164
rect 44 1172 400 1236
rect 44 762 108 1172
rect 400 1166 464 1172
rect 178 932 184 1100
rect 352 932 358 1100
rect 556 1096 748 1102
rect 184 658 352 932
rect 556 634 748 904
rect -1094 -44 -902 298
rect -1222 -108 436 -44
rect 500 -108 506 -44
rect -1222 -302 -1158 -108
rect -1094 -538 -902 -108
rect 556 -422 748 298
rect 814 -44 878 -38
rect 814 -282 878 -108
rect -1222 -1020 -1158 -690
rect -1222 -1110 -1158 -1084
rect -710 -1429 -524 -716
rect -460 -1084 -454 -1020
rect -390 -1084 -384 -1020
rect -454 -1262 -390 -1084
rect 38 -1134 44 -1070
rect 108 -1134 114 -1070
rect 44 -1278 108 -1134
rect 172 -1424 364 -758
rect 812 -1070 876 -894
rect 812 -1146 876 -1134
rect -1094 -2114 -902 -1726
rect -1094 -2294 -1088 -2114
rect -908 -2294 -902 -2114
rect -1094 -2306 -902 -2294
rect 556 -2110 748 -1726
rect 556 -2290 562 -2110
rect 742 -2290 748 -2110
rect 556 -2302 748 -2290
<< via1 >>
rect -454 1508 -390 1572
rect 44 1508 108 1572
rect -826 1164 -762 1228
rect -700 932 -532 1100
rect 400 1172 464 1236
rect 184 932 352 1100
rect 556 904 748 1096
rect 436 -108 500 -44
rect 814 -108 878 -44
rect -1222 -1084 -1158 -1020
rect -454 -1084 -390 -1020
rect 44 -1134 108 -1070
rect 812 -1134 876 -1070
<< metal2 >>
rect -826 1228 -762 2838
rect -454 1572 -390 1578
rect -390 1508 44 1572
rect 108 1508 114 1572
rect -454 1502 -390 1508
rect 400 1236 464 3056
rect -832 1164 -826 1228
rect -762 1164 -756 1228
rect 394 1172 400 1236
rect 464 1172 470 1236
rect 184 1100 352 1106
rect -706 932 -700 1100
rect -532 932 184 1100
rect 556 1096 748 2870
rect 184 926 352 932
rect 550 904 556 1096
rect 748 904 754 1096
rect 436 -44 500 -38
rect 500 -108 814 -44
rect 878 -108 884 -44
rect 436 -114 500 -108
rect -454 -1020 -390 -1014
rect -1228 -1084 -1222 -1020
rect -1158 -1084 -454 -1020
rect -454 -1090 -390 -1084
rect 44 -1070 108 -1064
rect 108 -1134 812 -1070
rect 876 -1134 882 -1070
rect 44 -1140 108 -1134
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ~/pro/aicex/ip/jnw_gr04_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1382 0 1 -990
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform -1 0 -230 0 1 -1958
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform -1 0 1036 0 1 -990
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 1 0 -116 0 1 -1958
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  JNWATR_PCH_4C1F2_0 ~/pro/aicex/ip/jnw_gr04_sky130a/design/JNW_ATR_SKY130A
timestamp 1744227008
transform 1 0 -116 0 1 66
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  JNWATR_PCH_4C1F2_1
timestamp 1744227008
transform -1 0 -230 0 1 66
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  JNWATR_PCH_4C1F2_2
timestamp 1744227008
transform -1 0 -230 0 1 1408
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  JNWATR_PCH_4C1F2_4
timestamp 1744227008
transform 1 0 -116 0 1 1408
box -184 -128 1336 928
use JNWTR_RPPO4  JNWTR_RPPO4_0 ~/pro/aicex/ip/jnw_gr04_sky130a/design/JNW_TR_SKY130A
timestamp 1744227008
transform -1 0 3248 0 1 -1642
box 0 0 1880 3440
<< labels >>
flabel locali -292 2488 -52 3066 0 FreeSans 1600 0 0 0 VDD
flabel locali 940 2850 1132 3042 0 FreeSans 1600 0 0 0 VSS
flabel metal2 556 2678 748 2870 0 FreeSans 1600 0 0 0 Vo
flabel metal2 400 2992 464 3056 0 FreeSans 1600 0 0 0 VIN
flabel metal2 -826 2768 -762 2832 0 FreeSans 1600 0 0 0 VIP
<< end >>
