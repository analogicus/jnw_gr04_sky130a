*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/PTAT_TO_COMP_lpe.spi
#else
.include ../../../work/xsch/PTAT_TO_COMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param vdda = 1.8
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc 1.8
V_I  OUT  0  dc  0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

* Translate names
VB0 temp.0 temp<0> dc 0
VB1 temp.1 temp<1> dc 0
VB2 temp.2 temp<2> dc 0
VB3 temp.3 temp<3> dc 0
VB4 temp.4 temp<4> dc 0
VB5 temp.5 temp<5> dc 0
VB6 temp.6 temp<6> dc 0
VB7 temp.7 temp<7> dc 0
VB8 comp_reset comp_reset<0> dc 0

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.option savecurrents
.save VD1_OUT
.save VD2_OUT

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control

set num_threads=8
set color0=white
set color1=black
unset askquit


*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low =te 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )


optran 0 0 0 1n 1u 0


set fend = .raw
foreach vtemp -40 -30 -20 -10 0 10 20 30 40 50 60 70 80 90 100 110 120
  option temp=$vtemp
  tran 1n 5u 10n
  write {cicname}_$vtemp$fend
end

quit

.endc

.end
