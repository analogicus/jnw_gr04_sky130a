magic
tech sky130A
magscale 1 2
timestamp 1744371203
<< locali >>
rect 5372 6244 5666 6273
rect 5372 6160 5440 6244
rect 4220 6088 5440 6160
rect 5596 6160 5666 6244
rect 5596 6088 6816 6160
rect 4220 5968 6816 6088
rect 4220 5808 4412 5968
rect 5372 5760 5666 5968
rect 2634 4728 2874 5218
rect 3962 5120 4074 5462
rect 4220 4502 4412 5360
rect 5372 5298 5612 5360
rect 5372 4474 5666 5298
rect 6626 4528 6818 5312
rect 5426 4450 5666 4474
rect 4220 1936 4412 2148
rect 3922 1824 4412 1936
rect 4220 1792 4412 1824
rect 5372 1792 5666 2196
rect 6626 1792 6818 2148
rect 4220 1786 6818 1792
rect 4220 1606 4994 1786
rect 5174 1606 5864 1786
rect 6044 1606 6818 1786
rect 4220 1600 6818 1606
<< viali >>
rect 5440 6088 5596 6244
rect 3518 4764 3698 4944
rect 4994 1606 5174 1786
rect 5864 1606 6044 1786
<< metal1 >>
rect 4992 6418 6026 6420
rect 4992 6252 6050 6418
rect 4992 5752 5160 6252
rect 5434 6244 5602 6252
rect 5434 6088 5440 6244
rect 5596 6088 5602 6244
rect 5434 6076 5602 6088
rect 5858 5752 6050 6252
rect 4604 5064 4796 5454
rect 5244 5064 5308 5296
rect 5730 5064 5794 5264
rect 4602 5000 5794 5064
rect 4604 4950 4796 5000
rect 3506 4944 4796 4950
rect 3506 4764 3518 4944
rect 3698 4764 4796 4944
rect 6242 4934 6434 5392
rect 5008 4932 6434 4934
rect 3506 4758 4796 4764
rect 5000 4766 6434 4932
rect 5000 4442 5168 4766
rect 5862 4630 6050 4766
rect 5858 4442 6050 4630
rect 4604 3714 4796 4058
rect 5244 3790 5308 3954
rect 5730 3786 5794 3954
rect 4604 3650 5794 3714
rect 4604 3334 4796 3650
rect 5244 3486 5308 3650
rect 5730 3490 5794 3650
rect 6242 3258 6434 4136
rect 4604 2564 4796 3088
rect 4988 2360 5180 3184
rect 5244 2686 5308 2894
rect 5730 2738 5794 2978
rect 5730 2642 5794 2732
rect 5858 2366 6050 3124
rect 6242 2484 6434 3026
rect 4988 1786 5180 2300
rect 4988 1606 4994 1786
rect 5174 1606 5180 1786
rect 4988 1594 5180 1606
rect 5858 1786 6050 2300
rect 5858 1606 5864 1786
rect 6044 1606 6050 1786
rect 5858 1594 6050 1606
use JNWTR_RPPO4  x2 ../JNW_TR_SKY130A
timestamp 1744227008
transform -1 0 4102 0 1 1808
box 0 0 1880 3440
use JNWATR_PCH_4C1F2  xb1 ../JNW_ATR_SKY130A
timestamp 1744227008
transform -1 0 5468 0 1 5160
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xb2
timestamp 1744227008
transform 1 0 5570 0 1 5160
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xi1
timestamp 1744227008
transform -1 0 5468 0 1 3850
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xi2
timestamp 1744227008
transform 1 0 5570 0 1 3850
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xm1_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform -1 0 5468 0 1 1996
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xm1_1
timestamp 1734044400
transform -1 0 5468 0 1 2794
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xm2_0
timestamp 1734044400
transform 1 0 5570 0 1 1996
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xm2_1
timestamp 1734044400
transform 1 0 5570 0 1 2794
box -184 -128 1336 928
<< labels >>
flabel metal1 5730 3786 5794 3954 0 FreeSans 1600 0 0 0 VIN
port 2 nsew
flabel metal1 5244 3790 5308 3954 0 FreeSans 1600 0 0 0 VIP
port 3 nsew
flabel metal1 6242 3258 6434 4136 0 FreeSans 1600 0 0 0 Vo
port 4 nsew
flabel metal1 4992 6252 5842 6420 0 FreeSans 1600 0 0 0 VDD
port 7 nsew
flabel metal1 5858 6220 6050 6412 0 FreeSans 1600 0 0 0 VDD
port 9 nsew
flabel locali 3962 5350 4074 5462 0 FreeSans 1600 0 0 0 VSS
port 11 nsew
<< end >>
