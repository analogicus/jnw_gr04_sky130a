magic
tech sky130A
timestamp 1743680127
<< end >>
